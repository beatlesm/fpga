module changevalue (
	output gps_lock
);

assign gps_lock = 1'b1;
endmodule
