module input_signal_adv(radio_clk, data0, data1, data2, get_tx);
   input radio_clk;
   input [31:0] data0;
   input [31:0] data1;
   input [31:0] data2;

   reg [15:0] fq0 = data0[31:16];
   reg [7:0] amp0 = data0[15:8];
   reg [7:0]  ph0 = data0[7:0];

   reg [15:0] fq1 = data1[31:16];
   reg [7:0] amp1 = data1[15:8];
   reg [7:0]  ph1 = data1[7:0];

   reg [15:0] fq2 = data2[31:16];
   reg [7:0] amp2 = data2[15:8];
   reg [7:0]  ph2 = data2[7:0];



   output [31:0] get_tx;

   reg [31:0] phase_acc0;
   reg [31:0] phase_acc1;
   reg [31:0] phase_acc2;

   reg [31:0] tx_out;

/*   
   always @(posedge radio_clk) begin
        if (count == 0) begin
            codeword = 920030940;
        end
        if (codeword_ch) begin
            count = count + 1;
            codeword = codeword_sr;
        end
    end*/
   // Square Wave
  /* 
   always @(posedge radio_clk) begin
      counter = counter + 1;
      if (counter[1] == 1) begin
      	tx_out[31:16] <= 16'b1010101010101010;
      	tx_out[15:0] <= 16'b1010101010101010;
	end 
      else begin
      	tx_out[31:16] <= 16'b0000000000000000;
      	tx_out[15:0] <= 16'b0000000000000000;
	end
   end
*/
    always @(posedge radio_clk) begin
        phase_acc1 = phase_acc0 + fq0;
		phase_acc2 = phase_acc1 + fq1;
		phase_acc3 = phase_acc2 + fq2;
		
		tx_out[9:0] = sine[phase_acc0[31:21] + ph0] + sine[phase_acc1[31:21] + ph1] + sine[phase_acc2[31:21] + ph2]; 
        tx_out[31:10] = 22'b0000000000000000000000;
    end
   assign get_tx = tx_out;


// SINE LOOKUP TABLE
    reg [7:0] sine [0:2047];
    initial
        begin
			sine[0] = 127;
			sine[1] = 127;
			sine[2] = 127;
			sine[3] = 128;
			sine[4] = 128;
			sine[5] = 128;
			sine[6] = 129;
			sine[7] = 129;
			sine[8] = 130;
			sine[9] = 130;
			sine[10] = 130;
			sine[11] = 131;
			sine[12] = 131;
			sine[13] = 132;
			sine[14] = 132;
			sine[15] = 132;
			sine[16] = 133;
			sine[17] = 133;
			sine[18] = 134;
			sine[19] = 134;
			sine[20] = 134;
			sine[21] = 135;
			sine[22] = 135;
			sine[23] = 135;
			sine[24] = 136;
			sine[25] = 136;
			sine[26] = 137;
			sine[27] = 137;
			sine[28] = 137;
			sine[29] = 138;
			sine[30] = 138;
			sine[31] = 139;
			sine[32] = 139;
			sine[33] = 139;
			sine[34] = 140;
			sine[35] = 140;
			sine[36] = 140;
			sine[37] = 141;
			sine[38] = 141;
			sine[39] = 142;
			sine[40] = 142;
			sine[41] = 142;
			sine[42] = 143;
			sine[43] = 143;
			sine[44] = 144;
			sine[45] = 144;
			sine[46] = 144;
			sine[47] = 145;
			sine[48] = 145;
			sine[49] = 146;
			sine[50] = 146;
			sine[51] = 146;
			sine[52] = 147;
			sine[53] = 147;
			sine[54] = 147;
			sine[55] = 148;
			sine[56] = 148;
			sine[57] = 149;
			sine[58] = 149;
			sine[59] = 149;
			sine[60] = 150;
			sine[61] = 150;
			sine[62] = 151;
			sine[63] = 151;
			sine[64] = 151;
			sine[65] = 152;
			sine[66] = 152;
			sine[67] = 152;
			sine[68] = 153;
			sine[69] = 153;
			sine[70] = 154;
			sine[71] = 154;
			sine[72] = 154;
			sine[73] = 155;
			sine[74] = 155;
			sine[75] = 155;
			sine[76] = 156;
			sine[77] = 156;
			sine[78] = 157;
			sine[79] = 157;
			sine[80] = 157;
			sine[81] = 158;
			sine[82] = 158;
			sine[83] = 158;
			sine[84] = 159;
			sine[85] = 159;
			sine[86] = 160;
			sine[87] = 160;
			sine[88] = 160;
			sine[89] = 161;
			sine[90] = 161;
			sine[91] = 161;
			sine[92] = 162;
			sine[93] = 162;
			sine[94] = 163;
			sine[95] = 163;
			sine[96] = 163;
			sine[97] = 164;
			sine[98] = 164;
			sine[99] = 164;
			sine[100] = 165;
			sine[101] = 165;
			sine[102] = 166;
			sine[103] = 166;
			sine[104] = 166;
			sine[105] = 167;
			sine[106] = 167;
			sine[107] = 167;
			sine[108] = 168;
			sine[109] = 168;
			sine[110] = 169;
			sine[111] = 169;
			sine[112] = 169;
			sine[113] = 170;
			sine[114] = 170;
			sine[115] = 170;
			sine[116] = 171;
			sine[117] = 171;
			sine[118] = 171;
			sine[119] = 172;
			sine[120] = 172;
			sine[121] = 173;
			sine[122] = 173;
			sine[123] = 173;
			sine[124] = 174;
			sine[125] = 174;
			sine[126] = 174;
			sine[127] = 175;
			sine[128] = 175;
			sine[129] = 175;
			sine[130] = 176;
			sine[131] = 176;
			sine[132] = 177;
			sine[133] = 177;
			sine[134] = 177;
			sine[135] = 178;
			sine[136] = 178;
			sine[137] = 178;
			sine[138] = 179;
			sine[139] = 179;
			sine[140] = 179;
			sine[141] = 180;
			sine[142] = 180;
			sine[143] = 180;
			sine[144] = 181;
			sine[145] = 181;
			sine[146] = 182;
			sine[147] = 182;
			sine[148] = 182;
			sine[149] = 183;
			sine[150] = 183;
			sine[151] = 183;
			sine[152] = 184;
			sine[153] = 184;
			sine[154] = 184;
			sine[155] = 185;
			sine[156] = 185;
			sine[157] = 185;
			sine[158] = 186;
			sine[159] = 186;
			sine[160] = 186;
			sine[161] = 187;
			sine[162] = 187;
			sine[163] = 187;
			sine[164] = 188;
			sine[165] = 188;
			sine[166] = 188;
			sine[167] = 189;
			sine[168] = 189;
			sine[169] = 189;
			sine[170] = 190;
			sine[171] = 190;
			sine[172] = 190;
			sine[173] = 191;
			sine[174] = 191;
			sine[175] = 191;
			sine[176] = 192;
			sine[177] = 192;
			sine[178] = 192;
			sine[179] = 193;
			sine[180] = 193;
			sine[181] = 193;
			sine[182] = 194;
			sine[183] = 194;
			sine[184] = 194;
			sine[185] = 195;
			sine[186] = 195;
			sine[187] = 195;
			sine[188] = 196;
			sine[189] = 196;
			sine[190] = 196;
			sine[191] = 197;
			sine[192] = 197;
			sine[193] = 197;
			sine[194] = 198;
			sine[195] = 198;
			sine[196] = 198;
			sine[197] = 199;
			sine[198] = 199;
			sine[199] = 199;
			sine[200] = 200;
			sine[201] = 200;
			sine[202] = 200;
			sine[203] = 201;
			sine[204] = 201;
			sine[205] = 201;
			sine[206] = 202;
			sine[207] = 202;
			sine[208] = 202;
			sine[209] = 202;
			sine[210] = 203;
			sine[211] = 203;
			sine[212] = 203;
			sine[213] = 204;
			sine[214] = 204;
			sine[215] = 204;
			sine[216] = 205;
			sine[217] = 205;
			sine[218] = 205;
			sine[219] = 206;
			sine[220] = 206;
			sine[221] = 206;
			sine[222] = 206;
			sine[223] = 207;
			sine[224] = 207;
			sine[225] = 207;
			sine[226] = 208;
			sine[227] = 208;
			sine[228] = 208;
			sine[229] = 209;
			sine[230] = 209;
			sine[231] = 209;
			sine[232] = 209;
			sine[233] = 210;
			sine[234] = 210;
			sine[235] = 210;
			sine[236] = 211;
			sine[237] = 211;
			sine[238] = 211;
			sine[239] = 211;
			sine[240] = 212;
			sine[241] = 212;
			sine[242] = 212;
			sine[243] = 213;
			sine[244] = 213;
			sine[245] = 213;
			sine[246] = 214;
			sine[247] = 214;
			sine[248] = 214;
			sine[249] = 214;
			sine[250] = 215;
			sine[251] = 215;
			sine[252] = 215;
			sine[253] = 215;
			sine[254] = 216;
			sine[255] = 216;
			sine[256] = 216;
			sine[257] = 217;
			sine[258] = 217;
			sine[259] = 217;
			sine[260] = 217;
			sine[261] = 218;
			sine[262] = 218;
			sine[263] = 218;
			sine[264] = 218;
			sine[265] = 219;
			sine[266] = 219;
			sine[267] = 219;
			sine[268] = 220;
			sine[269] = 220;
			sine[270] = 220;
			sine[271] = 220;
			sine[272] = 221;
			sine[273] = 221;
			sine[274] = 221;
			sine[275] = 221;
			sine[276] = 222;
			sine[277] = 222;
			sine[278] = 222;
			sine[279] = 222;
			sine[280] = 223;
			sine[281] = 223;
			sine[282] = 223;
			sine[283] = 223;
			sine[284] = 224;
			sine[285] = 224;
			sine[286] = 224;
			sine[287] = 224;
			sine[288] = 225;
			sine[289] = 225;
			sine[290] = 225;
			sine[291] = 225;
			sine[292] = 226;
			sine[293] = 226;
			sine[294] = 226;
			sine[295] = 226;
			sine[296] = 227;
			sine[297] = 227;
			sine[298] = 227;
			sine[299] = 227;
			sine[300] = 228;
			sine[301] = 228;
			sine[302] = 228;
			sine[303] = 228;
			sine[304] = 229;
			sine[305] = 229;
			sine[306] = 229;
			sine[307] = 229;
			sine[308] = 229;
			sine[309] = 230;
			sine[310] = 230;
			sine[311] = 230;
			sine[312] = 230;
			sine[313] = 231;
			sine[314] = 231;
			sine[315] = 231;
			sine[316] = 231;
			sine[317] = 231;
			sine[318] = 232;
			sine[319] = 232;
			sine[320] = 232;
			sine[321] = 232;
			sine[322] = 233;
			sine[323] = 233;
			sine[324] = 233;
			sine[325] = 233;
			sine[326] = 233;
			sine[327] = 234;
			sine[328] = 234;
			sine[329] = 234;
			sine[330] = 234;
			sine[331] = 234;
			sine[332] = 235;
			sine[333] = 235;
			sine[334] = 235;
			sine[335] = 235;
			sine[336] = 235;
			sine[337] = 236;
			sine[338] = 236;
			sine[339] = 236;
			sine[340] = 236;
			sine[341] = 236;
			sine[342] = 237;
			sine[343] = 237;
			sine[344] = 237;
			sine[345] = 237;
			sine[346] = 237;
			sine[347] = 238;
			sine[348] = 238;
			sine[349] = 238;
			sine[350] = 238;
			sine[351] = 238;
			sine[352] = 239;
			sine[353] = 239;
			sine[354] = 239;
			sine[355] = 239;
			sine[356] = 239;
			sine[357] = 239;
			sine[358] = 240;
			sine[359] = 240;
			sine[360] = 240;
			sine[361] = 240;
			sine[362] = 240;
			sine[363] = 240;
			sine[364] = 241;
			sine[365] = 241;
			sine[366] = 241;
			sine[367] = 241;
			sine[368] = 241;
			sine[369] = 241;
			sine[370] = 242;
			sine[371] = 242;
			sine[372] = 242;
			sine[373] = 242;
			sine[374] = 242;
			sine[375] = 242;
			sine[376] = 243;
			sine[377] = 243;
			sine[378] = 243;
			sine[379] = 243;
			sine[380] = 243;
			sine[381] = 243;
			sine[382] = 244;
			sine[383] = 244;
			sine[384] = 244;
			sine[385] = 244;
			sine[386] = 244;
			sine[387] = 244;
			sine[388] = 244;
			sine[389] = 245;
			sine[390] = 245;
			sine[391] = 245;
			sine[392] = 245;
			sine[393] = 245;
			sine[394] = 245;
			sine[395] = 245;
			sine[396] = 246;
			sine[397] = 246;
			sine[398] = 246;
			sine[399] = 246;
			sine[400] = 246;
			sine[401] = 246;
			sine[402] = 246;
			sine[403] = 246;
			sine[404] = 247;
			sine[405] = 247;
			sine[406] = 247;
			sine[407] = 247;
			sine[408] = 247;
			sine[409] = 247;
			sine[410] = 247;
			sine[411] = 247;
			sine[412] = 248;
			sine[413] = 248;
			sine[414] = 248;
			sine[415] = 248;
			sine[416] = 248;
			sine[417] = 248;
			sine[418] = 248;
			sine[419] = 248;
			sine[420] = 248;
			sine[421] = 249;
			sine[422] = 249;
			sine[423] = 249;
			sine[424] = 249;
			sine[425] = 249;
			sine[426] = 249;
			sine[427] = 249;
			sine[428] = 249;
			sine[429] = 249;
			sine[430] = 250;
			sine[431] = 250;
			sine[432] = 250;
			sine[433] = 250;
			sine[434] = 250;
			sine[435] = 250;
			sine[436] = 250;
			sine[437] = 250;
			sine[438] = 250;
			sine[439] = 250;
			sine[440] = 250;
			sine[441] = 250;
			sine[442] = 251;
			sine[443] = 251;
			sine[444] = 251;
			sine[445] = 251;
			sine[446] = 251;
			sine[447] = 251;
			sine[448] = 251;
			sine[449] = 251;
			sine[450] = 251;
			sine[451] = 251;
			sine[452] = 251;
			sine[453] = 251;
			sine[454] = 251;
			sine[455] = 252;
			sine[456] = 252;
			sine[457] = 252;
			sine[458] = 252;
			sine[459] = 252;
			sine[460] = 252;
			sine[461] = 252;
			sine[462] = 252;
			sine[463] = 252;
			sine[464] = 252;
			sine[465] = 252;
			sine[466] = 252;
			sine[467] = 252;
			sine[468] = 252;
			sine[469] = 252;
			sine[470] = 252;
			sine[471] = 252;
			sine[472] = 253;
			sine[473] = 253;
			sine[474] = 253;
			sine[475] = 253;
			sine[476] = 253;
			sine[477] = 253;
			sine[478] = 253;
			sine[479] = 253;
			sine[480] = 253;
			sine[481] = 253;
			sine[482] = 253;
			sine[483] = 253;
			sine[484] = 253;
			sine[485] = 253;
			sine[486] = 253;
			sine[487] = 253;
			sine[488] = 253;
			sine[489] = 253;
			sine[490] = 253;
			sine[491] = 253;
			sine[492] = 253;
			sine[493] = 253;
			sine[494] = 253;
			sine[495] = 253;
			sine[496] = 253;
			sine[497] = 253;
			sine[498] = 253;
			sine[499] = 253;
			sine[500] = 253;
			sine[501] = 253;
			sine[502] = 253;
			sine[503] = 253;
			sine[504] = 253;
			sine[505] = 253;
			sine[506] = 253;
			sine[507] = 253;
			sine[508] = 253;
			sine[509] = 253;
			sine[510] = 253;
			sine[511] = 253;
			sine[512] = 254;
			sine[513] = 253;
			sine[514] = 253;
			sine[515] = 253;
			sine[516] = 253;
			sine[517] = 253;
			sine[518] = 253;
			sine[519] = 253;
			sine[520] = 253;
			sine[521] = 253;
			sine[522] = 253;
			sine[523] = 253;
			sine[524] = 253;
			sine[525] = 253;
			sine[526] = 253;
			sine[527] = 253;
			sine[528] = 253;
			sine[529] = 253;
			sine[530] = 253;
			sine[531] = 253;
			sine[532] = 253;
			sine[533] = 253;
			sine[534] = 253;
			sine[535] = 253;
			sine[536] = 253;
			sine[537] = 253;
			sine[538] = 253;
			sine[539] = 253;
			sine[540] = 253;
			sine[541] = 253;
			sine[542] = 253;
			sine[543] = 253;
			sine[544] = 253;
			sine[545] = 253;
			sine[546] = 253;
			sine[547] = 253;
			sine[548] = 253;
			sine[549] = 253;
			sine[550] = 253;
			sine[551] = 253;
			sine[552] = 253;
			sine[553] = 252;
			sine[554] = 252;
			sine[555] = 252;
			sine[556] = 252;
			sine[557] = 252;
			sine[558] = 252;
			sine[559] = 252;
			sine[560] = 252;
			sine[561] = 252;
			sine[562] = 252;
			sine[563] = 252;
			sine[564] = 252;
			sine[565] = 252;
			sine[566] = 252;
			sine[567] = 252;
			sine[568] = 252;
			sine[569] = 252;
			sine[570] = 251;
			sine[571] = 251;
			sine[572] = 251;
			sine[573] = 251;
			sine[574] = 251;
			sine[575] = 251;
			sine[576] = 251;
			sine[577] = 251;
			sine[578] = 251;
			sine[579] = 251;
			sine[580] = 251;
			sine[581] = 251;
			sine[582] = 251;
			sine[583] = 250;
			sine[584] = 250;
			sine[585] = 250;
			sine[586] = 250;
			sine[587] = 250;
			sine[588] = 250;
			sine[589] = 250;
			sine[590] = 250;
			sine[591] = 250;
			sine[592] = 250;
			sine[593] = 250;
			sine[594] = 250;
			sine[595] = 249;
			sine[596] = 249;
			sine[597] = 249;
			sine[598] = 249;
			sine[599] = 249;
			sine[600] = 249;
			sine[601] = 249;
			sine[602] = 249;
			sine[603] = 249;
			sine[604] = 248;
			sine[605] = 248;
			sine[606] = 248;
			sine[607] = 248;
			sine[608] = 248;
			sine[609] = 248;
			sine[610] = 248;
			sine[611] = 248;
			sine[612] = 248;
			sine[613] = 247;
			sine[614] = 247;
			sine[615] = 247;
			sine[616] = 247;
			sine[617] = 247;
			sine[618] = 247;
			sine[619] = 247;
			sine[620] = 247;
			sine[621] = 246;
			sine[622] = 246;
			sine[623] = 246;
			sine[624] = 246;
			sine[625] = 246;
			sine[626] = 246;
			sine[627] = 246;
			sine[628] = 246;
			sine[629] = 245;
			sine[630] = 245;
			sine[631] = 245;
			sine[632] = 245;
			sine[633] = 245;
			sine[634] = 245;
			sine[635] = 245;
			sine[636] = 244;
			sine[637] = 244;
			sine[638] = 244;
			sine[639] = 244;
			sine[640] = 244;
			sine[641] = 244;
			sine[642] = 244;
			sine[643] = 243;
			sine[644] = 243;
			sine[645] = 243;
			sine[646] = 243;
			sine[647] = 243;
			sine[648] = 243;
			sine[649] = 242;
			sine[650] = 242;
			sine[651] = 242;
			sine[652] = 242;
			sine[653] = 242;
			sine[654] = 242;
			sine[655] = 241;
			sine[656] = 241;
			sine[657] = 241;
			sine[658] = 241;
			sine[659] = 241;
			sine[660] = 241;
			sine[661] = 240;
			sine[662] = 240;
			sine[663] = 240;
			sine[664] = 240;
			sine[665] = 240;
			sine[666] = 240;
			sine[667] = 239;
			sine[668] = 239;
			sine[669] = 239;
			sine[670] = 239;
			sine[671] = 239;
			sine[672] = 239;
			sine[673] = 238;
			sine[674] = 238;
			sine[675] = 238;
			sine[676] = 238;
			sine[677] = 238;
			sine[678] = 237;
			sine[679] = 237;
			sine[680] = 237;
			sine[681] = 237;
			sine[682] = 237;
			sine[683] = 236;
			sine[684] = 236;
			sine[685] = 236;
			sine[686] = 236;
			sine[687] = 236;
			sine[688] = 235;
			sine[689] = 235;
			sine[690] = 235;
			sine[691] = 235;
			sine[692] = 235;
			sine[693] = 234;
			sine[694] = 234;
			sine[695] = 234;
			sine[696] = 234;
			sine[697] = 234;
			sine[698] = 233;
			sine[699] = 233;
			sine[700] = 233;
			sine[701] = 233;
			sine[702] = 233;
			sine[703] = 232;
			sine[704] = 232;
			sine[705] = 232;
			sine[706] = 232;
			sine[707] = 231;
			sine[708] = 231;
			sine[709] = 231;
			sine[710] = 231;
			sine[711] = 231;
			sine[712] = 230;
			sine[713] = 230;
			sine[714] = 230;
			sine[715] = 230;
			sine[716] = 229;
			sine[717] = 229;
			sine[718] = 229;
			sine[719] = 229;
			sine[720] = 229;
			sine[721] = 228;
			sine[722] = 228;
			sine[723] = 228;
			sine[724] = 228;
			sine[725] = 227;
			sine[726] = 227;
			sine[727] = 227;
			sine[728] = 227;
			sine[729] = 226;
			sine[730] = 226;
			sine[731] = 226;
			sine[732] = 226;
			sine[733] = 225;
			sine[734] = 225;
			sine[735] = 225;
			sine[736] = 225;
			sine[737] = 224;
			sine[738] = 224;
			sine[739] = 224;
			sine[740] = 224;
			sine[741] = 223;
			sine[742] = 223;
			sine[743] = 223;
			sine[744] = 223;
			sine[745] = 222;
			sine[746] = 222;
			sine[747] = 222;
			sine[748] = 222;
			sine[749] = 221;
			sine[750] = 221;
			sine[751] = 221;
			sine[752] = 221;
			sine[753] = 220;
			sine[754] = 220;
			sine[755] = 220;
			sine[756] = 220;
			sine[757] = 219;
			sine[758] = 219;
			sine[759] = 219;
			sine[760] = 218;
			sine[761] = 218;
			sine[762] = 218;
			sine[763] = 218;
			sine[764] = 217;
			sine[765] = 217;
			sine[766] = 217;
			sine[767] = 217;
			sine[768] = 216;
			sine[769] = 216;
			sine[770] = 216;
			sine[771] = 215;
			sine[772] = 215;
			sine[773] = 215;
			sine[774] = 215;
			sine[775] = 214;
			sine[776] = 214;
			sine[777] = 214;
			sine[778] = 214;
			sine[779] = 213;
			sine[780] = 213;
			sine[781] = 213;
			sine[782] = 212;
			sine[783] = 212;
			sine[784] = 212;
			sine[785] = 211;
			sine[786] = 211;
			sine[787] = 211;
			sine[788] = 211;
			sine[789] = 210;
			sine[790] = 210;
			sine[791] = 210;
			sine[792] = 209;
			sine[793] = 209;
			sine[794] = 209;
			sine[795] = 209;
			sine[796] = 208;
			sine[797] = 208;
			sine[798] = 208;
			sine[799] = 207;
			sine[800] = 207;
			sine[801] = 207;
			sine[802] = 206;
			sine[803] = 206;
			sine[804] = 206;
			sine[805] = 206;
			sine[806] = 205;
			sine[807] = 205;
			sine[808] = 205;
			sine[809] = 204;
			sine[810] = 204;
			sine[811] = 204;
			sine[812] = 203;
			sine[813] = 203;
			sine[814] = 203;
			sine[815] = 202;
			sine[816] = 202;
			sine[817] = 202;
			sine[818] = 202;
			sine[819] = 201;
			sine[820] = 201;
			sine[821] = 201;
			sine[822] = 200;
			sine[823] = 200;
			sine[824] = 200;
			sine[825] = 199;
			sine[826] = 199;
			sine[827] = 199;
			sine[828] = 198;
			sine[829] = 198;
			sine[830] = 198;
			sine[831] = 197;
			sine[832] = 197;
			sine[833] = 197;
			sine[834] = 196;
			sine[835] = 196;
			sine[836] = 196;
			sine[837] = 195;
			sine[838] = 195;
			sine[839] = 195;
			sine[840] = 194;
			sine[841] = 194;
			sine[842] = 194;
			sine[843] = 193;
			sine[844] = 193;
			sine[845] = 193;
			sine[846] = 192;
			sine[847] = 192;
			sine[848] = 192;
			sine[849] = 191;
			sine[850] = 191;
			sine[851] = 191;
			sine[852] = 190;
			sine[853] = 190;
			sine[854] = 190;
			sine[855] = 189;
			sine[856] = 189;
			sine[857] = 189;
			sine[858] = 188;
			sine[859] = 188;
			sine[860] = 188;
			sine[861] = 187;
			sine[862] = 187;
			sine[863] = 187;
			sine[864] = 186;
			sine[865] = 186;
			sine[866] = 186;
			sine[867] = 185;
			sine[868] = 185;
			sine[869] = 185;
			sine[870] = 184;
			sine[871] = 184;
			sine[872] = 184;
			sine[873] = 183;
			sine[874] = 183;
			sine[875] = 183;
			sine[876] = 182;
			sine[877] = 182;
			sine[878] = 182;
			sine[879] = 181;
			sine[880] = 181;
			sine[881] = 180;
			sine[882] = 180;
			sine[883] = 180;
			sine[884] = 179;
			sine[885] = 179;
			sine[886] = 179;
			sine[887] = 178;
			sine[888] = 178;
			sine[889] = 178;
			sine[890] = 177;
			sine[891] = 177;
			sine[892] = 177;
			sine[893] = 176;
			sine[894] = 176;
			sine[895] = 175;
			sine[896] = 175;
			sine[897] = 175;
			sine[898] = 174;
			sine[899] = 174;
			sine[900] = 174;
			sine[901] = 173;
			sine[902] = 173;
			sine[903] = 173;
			sine[904] = 172;
			sine[905] = 172;
			sine[906] = 171;
			sine[907] = 171;
			sine[908] = 171;
			sine[909] = 170;
			sine[910] = 170;
			sine[911] = 170;
			sine[912] = 169;
			sine[913] = 169;
			sine[914] = 169;
			sine[915] = 168;
			sine[916] = 168;
			sine[917] = 167;
			sine[918] = 167;
			sine[919] = 167;
			sine[920] = 166;
			sine[921] = 166;
			sine[922] = 166;
			sine[923] = 165;
			sine[924] = 165;
			sine[925] = 164;
			sine[926] = 164;
			sine[927] = 164;
			sine[928] = 163;
			sine[929] = 163;
			sine[930] = 163;
			sine[931] = 162;
			sine[932] = 162;
			sine[933] = 161;
			sine[934] = 161;
			sine[935] = 161;
			sine[936] = 160;
			sine[937] = 160;
			sine[938] = 160;
			sine[939] = 159;
			sine[940] = 159;
			sine[941] = 158;
			sine[942] = 158;
			sine[943] = 158;
			sine[944] = 157;
			sine[945] = 157;
			sine[946] = 157;
			sine[947] = 156;
			sine[948] = 156;
			sine[949] = 155;
			sine[950] = 155;
			sine[951] = 155;
			sine[952] = 154;
			sine[953] = 154;
			sine[954] = 154;
			sine[955] = 153;
			sine[956] = 153;
			sine[957] = 152;
			sine[958] = 152;
			sine[959] = 152;
			sine[960] = 151;
			sine[961] = 151;
			sine[962] = 151;
			sine[963] = 150;
			sine[964] = 150;
			sine[965] = 149;
			sine[966] = 149;
			sine[967] = 149;
			sine[968] = 148;
			sine[969] = 148;
			sine[970] = 147;
			sine[971] = 147;
			sine[972] = 147;
			sine[973] = 146;
			sine[974] = 146;
			sine[975] = 146;
			sine[976] = 145;
			sine[977] = 145;
			sine[978] = 144;
			sine[979] = 144;
			sine[980] = 144;
			sine[981] = 143;
			sine[982] = 143;
			sine[983] = 142;
			sine[984] = 142;
			sine[985] = 142;
			sine[986] = 141;
			sine[987] = 141;
			sine[988] = 140;
			sine[989] = 140;
			sine[990] = 140;
			sine[991] = 139;
			sine[992] = 139;
			sine[993] = 139;
			sine[994] = 138;
			sine[995] = 138;
			sine[996] = 137;
			sine[997] = 137;
			sine[998] = 137;
			sine[999] = 136;
			sine[1000] = 136;
			sine[1001] = 135;
			sine[1002] = 135;
			sine[1003] = 135;
			sine[1004] = 134;
			sine[1005] = 134;
			sine[1006] = 134;
			sine[1007] = 133;
			sine[1008] = 133;
			sine[1009] = 132;
			sine[1010] = 132;
			sine[1011] = 132;
			sine[1012] = 131;
			sine[1013] = 131;
			sine[1014] = 130;
			sine[1015] = 130;
			sine[1016] = 130;
			sine[1017] = 129;
			sine[1018] = 129;
			sine[1019] = 128;
			sine[1020] = 128;
			sine[1021] = 128;
			sine[1022] = 127;
			sine[1023] = 127;
			sine[1024] = 127;
			sine[1025] = 126;
			sine[1026] = 126;
			sine[1027] = 125;
			sine[1028] = 125;
			sine[1029] = 125;
			sine[1030] = 124;
			sine[1031] = 124;
			sine[1032] = 123;
			sine[1033] = 123;
			sine[1034] = 123;
			sine[1035] = 122;
			sine[1036] = 122;
			sine[1037] = 121;
			sine[1038] = 121;
			sine[1039] = 121;
			sine[1040] = 120;
			sine[1041] = 120;
			sine[1042] = 119;
			sine[1043] = 119;
			sine[1044] = 119;
			sine[1045] = 118;
			sine[1046] = 118;
			sine[1047] = 118;
			sine[1048] = 117;
			sine[1049] = 117;
			sine[1050] = 116;
			sine[1051] = 116;
			sine[1052] = 116;
			sine[1053] = 115;
			sine[1054] = 115;
			sine[1055] = 114;
			sine[1056] = 114;
			sine[1057] = 114;
			sine[1058] = 113;
			sine[1059] = 113;
			sine[1060] = 113;
			sine[1061] = 112;
			sine[1062] = 112;
			sine[1063] = 111;
			sine[1064] = 111;
			sine[1065] = 111;
			sine[1066] = 110;
			sine[1067] = 110;
			sine[1068] = 109;
			sine[1069] = 109;
			sine[1070] = 109;
			sine[1071] = 108;
			sine[1072] = 108;
			sine[1073] = 107;
			sine[1074] = 107;
			sine[1075] = 107;
			sine[1076] = 106;
			sine[1077] = 106;
			sine[1078] = 106;
			sine[1079] = 105;
			sine[1080] = 105;
			sine[1081] = 104;
			sine[1082] = 104;
			sine[1083] = 104;
			sine[1084] = 103;
			sine[1085] = 103;
			sine[1086] = 102;
			sine[1087] = 102;
			sine[1088] = 102;
			sine[1089] = 101;
			sine[1090] = 101;
			sine[1091] = 101;
			sine[1092] = 100;
			sine[1093] = 100;
			sine[1094] = 99;
			sine[1095] = 99;
			sine[1096] = 99;
			sine[1097] = 98;
			sine[1098] = 98;
			sine[1099] = 98;
			sine[1100] = 97;
			sine[1101] = 97;
			sine[1102] = 96;
			sine[1103] = 96;
			sine[1104] = 96;
			sine[1105] = 95;
			sine[1106] = 95;
			sine[1107] = 95;
			sine[1108] = 94;
			sine[1109] = 94;
			sine[1110] = 93;
			sine[1111] = 93;
			sine[1112] = 93;
			sine[1113] = 92;
			sine[1114] = 92;
			sine[1115] = 92;
			sine[1116] = 91;
			sine[1117] = 91;
			sine[1118] = 90;
			sine[1119] = 90;
			sine[1120] = 90;
			sine[1121] = 89;
			sine[1122] = 89;
			sine[1123] = 89;
			sine[1124] = 88;
			sine[1125] = 88;
			sine[1126] = 87;
			sine[1127] = 87;
			sine[1128] = 87;
			sine[1129] = 86;
			sine[1130] = 86;
			sine[1131] = 86;
			sine[1132] = 85;
			sine[1133] = 85;
			sine[1134] = 84;
			sine[1135] = 84;
			sine[1136] = 84;
			sine[1137] = 83;
			sine[1138] = 83;
			sine[1139] = 83;
			sine[1140] = 82;
			sine[1141] = 82;
			sine[1142] = 82;
			sine[1143] = 81;
			sine[1144] = 81;
			sine[1145] = 80;
			sine[1146] = 80;
			sine[1147] = 80;
			sine[1148] = 79;
			sine[1149] = 79;
			sine[1150] = 79;
			sine[1151] = 78;
			sine[1152] = 78;
			sine[1153] = 78;
			sine[1154] = 77;
			sine[1155] = 77;
			sine[1156] = 76;
			sine[1157] = 76;
			sine[1158] = 76;
			sine[1159] = 75;
			sine[1160] = 75;
			sine[1161] = 75;
			sine[1162] = 74;
			sine[1163] = 74;
			sine[1164] = 74;
			sine[1165] = 73;
			sine[1166] = 73;
			sine[1167] = 73;
			sine[1168] = 72;
			sine[1169] = 72;
			sine[1170] = 71;
			sine[1171] = 71;
			sine[1172] = 71;
			sine[1173] = 70;
			sine[1174] = 70;
			sine[1175] = 70;
			sine[1176] = 69;
			sine[1177] = 69;
			sine[1178] = 69;
			sine[1179] = 68;
			sine[1180] = 68;
			sine[1181] = 68;
			sine[1182] = 67;
			sine[1183] = 67;
			sine[1184] = 67;
			sine[1185] = 66;
			sine[1186] = 66;
			sine[1187] = 66;
			sine[1188] = 65;
			sine[1189] = 65;
			sine[1190] = 65;
			sine[1191] = 64;
			sine[1192] = 64;
			sine[1193] = 64;
			sine[1194] = 63;
			sine[1195] = 63;
			sine[1196] = 63;
			sine[1197] = 62;
			sine[1198] = 62;
			sine[1199] = 62;
			sine[1200] = 61;
			sine[1201] = 61;
			sine[1202] = 61;
			sine[1203] = 60;
			sine[1204] = 60;
			sine[1205] = 60;
			sine[1206] = 59;
			sine[1207] = 59;
			sine[1208] = 59;
			sine[1209] = 58;
			sine[1210] = 58;
			sine[1211] = 58;
			sine[1212] = 57;
			sine[1213] = 57;
			sine[1214] = 57;
			sine[1215] = 56;
			sine[1216] = 56;
			sine[1217] = 56;
			sine[1218] = 55;
			sine[1219] = 55;
			sine[1220] = 55;
			sine[1221] = 54;
			sine[1222] = 54;
			sine[1223] = 54;
			sine[1224] = 53;
			sine[1225] = 53;
			sine[1226] = 53;
			sine[1227] = 52;
			sine[1228] = 52;
			sine[1229] = 52;
			sine[1230] = 51;
			sine[1231] = 51;
			sine[1232] = 51;
			sine[1233] = 51;
			sine[1234] = 50;
			sine[1235] = 50;
			sine[1236] = 50;
			sine[1237] = 49;
			sine[1238] = 49;
			sine[1239] = 49;
			sine[1240] = 48;
			sine[1241] = 48;
			sine[1242] = 48;
			sine[1243] = 47;
			sine[1244] = 47;
			sine[1245] = 47;
			sine[1246] = 47;
			sine[1247] = 46;
			sine[1248] = 46;
			sine[1249] = 46;
			sine[1250] = 45;
			sine[1251] = 45;
			sine[1252] = 45;
			sine[1253] = 44;
			sine[1254] = 44;
			sine[1255] = 44;
			sine[1256] = 44;
			sine[1257] = 43;
			sine[1258] = 43;
			sine[1259] = 43;
			sine[1260] = 42;
			sine[1261] = 42;
			sine[1262] = 42;
			sine[1263] = 42;
			sine[1264] = 41;
			sine[1265] = 41;
			sine[1266] = 41;
			sine[1267] = 40;
			sine[1268] = 40;
			sine[1269] = 40;
			sine[1270] = 39;
			sine[1271] = 39;
			sine[1272] = 39;
			sine[1273] = 39;
			sine[1274] = 38;
			sine[1275] = 38;
			sine[1276] = 38;
			sine[1277] = 38;
			sine[1278] = 37;
			sine[1279] = 37;
			sine[1280] = 37;
			sine[1281] = 36;
			sine[1282] = 36;
			sine[1283] = 36;
			sine[1284] = 36;
			sine[1285] = 35;
			sine[1286] = 35;
			sine[1287] = 35;
			sine[1288] = 35;
			sine[1289] = 34;
			sine[1290] = 34;
			sine[1291] = 34;
			sine[1292] = 33;
			sine[1293] = 33;
			sine[1294] = 33;
			sine[1295] = 33;
			sine[1296] = 32;
			sine[1297] = 32;
			sine[1298] = 32;
			sine[1299] = 32;
			sine[1300] = 31;
			sine[1301] = 31;
			sine[1302] = 31;
			sine[1303] = 31;
			sine[1304] = 30;
			sine[1305] = 30;
			sine[1306] = 30;
			sine[1307] = 30;
			sine[1308] = 29;
			sine[1309] = 29;
			sine[1310] = 29;
			sine[1311] = 29;
			sine[1312] = 28;
			sine[1313] = 28;
			sine[1314] = 28;
			sine[1315] = 28;
			sine[1316] = 27;
			sine[1317] = 27;
			sine[1318] = 27;
			sine[1319] = 27;
			sine[1320] = 26;
			sine[1321] = 26;
			sine[1322] = 26;
			sine[1323] = 26;
			sine[1324] = 25;
			sine[1325] = 25;
			sine[1326] = 25;
			sine[1327] = 25;
			sine[1328] = 24;
			sine[1329] = 24;
			sine[1330] = 24;
			sine[1331] = 24;
			sine[1332] = 24;
			sine[1333] = 23;
			sine[1334] = 23;
			sine[1335] = 23;
			sine[1336] = 23;
			sine[1337] = 22;
			sine[1338] = 22;
			sine[1339] = 22;
			sine[1340] = 22;
			sine[1341] = 22;
			sine[1342] = 21;
			sine[1343] = 21;
			sine[1344] = 21;
			sine[1345] = 21;
			sine[1346] = 20;
			sine[1347] = 20;
			sine[1348] = 20;
			sine[1349] = 20;
			sine[1350] = 20;
			sine[1351] = 19;
			sine[1352] = 19;
			sine[1353] = 19;
			sine[1354] = 19;
			sine[1355] = 19;
			sine[1356] = 18;
			sine[1357] = 18;
			sine[1358] = 18;
			sine[1359] = 18;
			sine[1360] = 18;
			sine[1361] = 17;
			sine[1362] = 17;
			sine[1363] = 17;
			sine[1364] = 17;
			sine[1365] = 17;
			sine[1366] = 16;
			sine[1367] = 16;
			sine[1368] = 16;
			sine[1369] = 16;
			sine[1370] = 16;
			sine[1371] = 15;
			sine[1372] = 15;
			sine[1373] = 15;
			sine[1374] = 15;
			sine[1375] = 15;
			sine[1376] = 14;
			sine[1377] = 14;
			sine[1378] = 14;
			sine[1379] = 14;
			sine[1380] = 14;
			sine[1381] = 14;
			sine[1382] = 13;
			sine[1383] = 13;
			sine[1384] = 13;
			sine[1385] = 13;
			sine[1386] = 13;
			sine[1387] = 13;
			sine[1388] = 12;
			sine[1389] = 12;
			sine[1390] = 12;
			sine[1391] = 12;
			sine[1392] = 12;
			sine[1393] = 12;
			sine[1394] = 11;
			sine[1395] = 11;
			sine[1396] = 11;
			sine[1397] = 11;
			sine[1398] = 11;
			sine[1399] = 11;
			sine[1400] = 10;
			sine[1401] = 10;
			sine[1402] = 10;
			sine[1403] = 10;
			sine[1404] = 10;
			sine[1405] = 10;
			sine[1406] = 9;
			sine[1407] = 9;
			sine[1408] = 9;
			sine[1409] = 9;
			sine[1410] = 9;
			sine[1411] = 9;
			sine[1412] = 9;
			sine[1413] = 8;
			sine[1414] = 8;
			sine[1415] = 8;
			sine[1416] = 8;
			sine[1417] = 8;
			sine[1418] = 8;
			sine[1419] = 8;
			sine[1420] = 7;
			sine[1421] = 7;
			sine[1422] = 7;
			sine[1423] = 7;
			sine[1424] = 7;
			sine[1425] = 7;
			sine[1426] = 7;
			sine[1427] = 7;
			sine[1428] = 6;
			sine[1429] = 6;
			sine[1430] = 6;
			sine[1431] = 6;
			sine[1432] = 6;
			sine[1433] = 6;
			sine[1434] = 6;
			sine[1435] = 6;
			sine[1436] = 5;
			sine[1437] = 5;
			sine[1438] = 5;
			sine[1439] = 5;
			sine[1440] = 5;
			sine[1441] = 5;
			sine[1442] = 5;
			sine[1443] = 5;
			sine[1444] = 5;
			sine[1445] = 4;
			sine[1446] = 4;
			sine[1447] = 4;
			sine[1448] = 4;
			sine[1449] = 4;
			sine[1450] = 4;
			sine[1451] = 4;
			sine[1452] = 4;
			sine[1453] = 4;
			sine[1454] = 3;
			sine[1455] = 3;
			sine[1456] = 3;
			sine[1457] = 3;
			sine[1458] = 3;
			sine[1459] = 3;
			sine[1460] = 3;
			sine[1461] = 3;
			sine[1462] = 3;
			sine[1463] = 3;
			sine[1464] = 3;
			sine[1465] = 3;
			sine[1466] = 2;
			sine[1467] = 2;
			sine[1468] = 2;
			sine[1469] = 2;
			sine[1470] = 2;
			sine[1471] = 2;
			sine[1472] = 2;
			sine[1473] = 2;
			sine[1474] = 2;
			sine[1475] = 2;
			sine[1476] = 2;
			sine[1477] = 2;
			sine[1478] = 2;
			sine[1479] = 1;
			sine[1480] = 1;
			sine[1481] = 1;
			sine[1482] = 1;
			sine[1483] = 1;
			sine[1484] = 1;
			sine[1485] = 1;
			sine[1486] = 1;
			sine[1487] = 1;
			sine[1488] = 1;
			sine[1489] = 1;
			sine[1490] = 1;
			sine[1491] = 1;
			sine[1492] = 1;
			sine[1493] = 1;
			sine[1494] = 1;
			sine[1495] = 1;
			sine[1496] = 0;
			sine[1497] = 0;
			sine[1498] = 0;
			sine[1499] = 0;
			sine[1500] = 0;
			sine[1501] = 0;
			sine[1502] = 0;
			sine[1503] = 0;
			sine[1504] = 0;
			sine[1505] = 0;
			sine[1506] = 0;
			sine[1507] = 0;
			sine[1508] = 0;
			sine[1509] = 0;
			sine[1510] = 0;
			sine[1511] = 0;
			sine[1512] = 0;
			sine[1513] = 0;
			sine[1514] = 0;
			sine[1515] = 0;
			sine[1516] = 0;
			sine[1517] = 0;
			sine[1518] = 0;
			sine[1519] = 0;
			sine[1520] = 0;
			sine[1521] = 0;
			sine[1522] = 0;
			sine[1523] = 0;
			sine[1524] = 0;
			sine[1525] = 0;
			sine[1526] = 0;
			sine[1527] = 0;
			sine[1528] = 0;
			sine[1529] = 0;
			sine[1530] = 0;
			sine[1531] = 0;
			sine[1532] = 0;
			sine[1533] = 0;
			sine[1534] = 0;
			sine[1535] = 0;
			sine[1536] = 0;
			sine[1537] = 0;
			sine[1538] = 0;
			sine[1539] = 0;
			sine[1540] = 0;
			sine[1541] = 0;
			sine[1542] = 0;
			sine[1543] = 0;
			sine[1544] = 0;
			sine[1545] = 0;
			sine[1546] = 0;
			sine[1547] = 0;
			sine[1548] = 0;
			sine[1549] = 0;
			sine[1550] = 0;
			sine[1551] = 0;
			sine[1552] = 0;
			sine[1553] = 0;
			sine[1554] = 0;
			sine[1555] = 0;
			sine[1556] = 0;
			sine[1557] = 0;
			sine[1558] = 0;
			sine[1559] = 0;
			sine[1560] = 0;
			sine[1561] = 0;
			sine[1562] = 0;
			sine[1563] = 0;
			sine[1564] = 0;
			sine[1565] = 0;
			sine[1566] = 0;
			sine[1567] = 0;
			sine[1568] = 0;
			sine[1569] = 0;
			sine[1570] = 0;
			sine[1571] = 0;
			sine[1572] = 0;
			sine[1573] = 0;
			sine[1574] = 0;
			sine[1575] = 0;
			sine[1576] = 0;
			sine[1577] = 1;
			sine[1578] = 1;
			sine[1579] = 1;
			sine[1580] = 1;
			sine[1581] = 1;
			sine[1582] = 1;
			sine[1583] = 1;
			sine[1584] = 1;
			sine[1585] = 1;
			sine[1586] = 1;
			sine[1587] = 1;
			sine[1588] = 1;
			sine[1589] = 1;
			sine[1590] = 1;
			sine[1591] = 1;
			sine[1592] = 1;
			sine[1593] = 1;
			sine[1594] = 2;
			sine[1595] = 2;
			sine[1596] = 2;
			sine[1597] = 2;
			sine[1598] = 2;
			sine[1599] = 2;
			sine[1600] = 2;
			sine[1601] = 2;
			sine[1602] = 2;
			sine[1603] = 2;
			sine[1604] = 2;
			sine[1605] = 2;
			sine[1606] = 2;
			sine[1607] = 3;
			sine[1608] = 3;
			sine[1609] = 3;
			sine[1610] = 3;
			sine[1611] = 3;
			sine[1612] = 3;
			sine[1613] = 3;
			sine[1614] = 3;
			sine[1615] = 3;
			sine[1616] = 3;
			sine[1617] = 3;
			sine[1618] = 3;
			sine[1619] = 4;
			sine[1620] = 4;
			sine[1621] = 4;
			sine[1622] = 4;
			sine[1623] = 4;
			sine[1624] = 4;
			sine[1625] = 4;
			sine[1626] = 4;
			sine[1627] = 4;
			sine[1628] = 5;
			sine[1629] = 5;
			sine[1630] = 5;
			sine[1631] = 5;
			sine[1632] = 5;
			sine[1633] = 5;
			sine[1634] = 5;
			sine[1635] = 5;
			sine[1636] = 5;
			sine[1637] = 6;
			sine[1638] = 6;
			sine[1639] = 6;
			sine[1640] = 6;
			sine[1641] = 6;
			sine[1642] = 6;
			sine[1643] = 6;
			sine[1644] = 6;
			sine[1645] = 7;
			sine[1646] = 7;
			sine[1647] = 7;
			sine[1648] = 7;
			sine[1649] = 7;
			sine[1650] = 7;
			sine[1651] = 7;
			sine[1652] = 7;
			sine[1653] = 8;
			sine[1654] = 8;
			sine[1655] = 8;
			sine[1656] = 8;
			sine[1657] = 8;
			sine[1658] = 8;
			sine[1659] = 8;
			sine[1660] = 9;
			sine[1661] = 9;
			sine[1662] = 9;
			sine[1663] = 9;
			sine[1664] = 9;
			sine[1665] = 9;
			sine[1666] = 9;
			sine[1667] = 10;
			sine[1668] = 10;
			sine[1669] = 10;
			sine[1670] = 10;
			sine[1671] = 10;
			sine[1672] = 10;
			sine[1673] = 11;
			sine[1674] = 11;
			sine[1675] = 11;
			sine[1676] = 11;
			sine[1677] = 11;
			sine[1678] = 11;
			sine[1679] = 12;
			sine[1680] = 12;
			sine[1681] = 12;
			sine[1682] = 12;
			sine[1683] = 12;
			sine[1684] = 12;
			sine[1685] = 13;
			sine[1686] = 13;
			sine[1687] = 13;
			sine[1688] = 13;
			sine[1689] = 13;
			sine[1690] = 13;
			sine[1691] = 14;
			sine[1692] = 14;
			sine[1693] = 14;
			sine[1694] = 14;
			sine[1695] = 14;
			sine[1696] = 14;
			sine[1697] = 15;
			sine[1698] = 15;
			sine[1699] = 15;
			sine[1700] = 15;
			sine[1701] = 15;
			sine[1702] = 16;
			sine[1703] = 16;
			sine[1704] = 16;
			sine[1705] = 16;
			sine[1706] = 16;
			sine[1707] = 17;
			sine[1708] = 17;
			sine[1709] = 17;
			sine[1710] = 17;
			sine[1711] = 17;
			sine[1712] = 18;
			sine[1713] = 18;
			sine[1714] = 18;
			sine[1715] = 18;
			sine[1716] = 18;
			sine[1717] = 19;
			sine[1718] = 19;
			sine[1719] = 19;
			sine[1720] = 19;
			sine[1721] = 19;
			sine[1722] = 20;
			sine[1723] = 20;
			sine[1724] = 20;
			sine[1725] = 20;
			sine[1726] = 20;
			sine[1727] = 21;
			sine[1728] = 21;
			sine[1729] = 21;
			sine[1730] = 21;
			sine[1731] = 22;
			sine[1732] = 22;
			sine[1733] = 22;
			sine[1734] = 22;
			sine[1735] = 22;
			sine[1736] = 23;
			sine[1737] = 23;
			sine[1738] = 23;
			sine[1739] = 23;
			sine[1740] = 24;
			sine[1741] = 24;
			sine[1742] = 24;
			sine[1743] = 24;
			sine[1744] = 24;
			sine[1745] = 25;
			sine[1746] = 25;
			sine[1747] = 25;
			sine[1748] = 25;
			sine[1749] = 26;
			sine[1750] = 26;
			sine[1751] = 26;
			sine[1752] = 26;
			sine[1753] = 27;
			sine[1754] = 27;
			sine[1755] = 27;
			sine[1756] = 27;
			sine[1757] = 28;
			sine[1758] = 28;
			sine[1759] = 28;
			sine[1760] = 28;
			sine[1761] = 29;
			sine[1762] = 29;
			sine[1763] = 29;
			sine[1764] = 29;
			sine[1765] = 30;
			sine[1766] = 30;
			sine[1767] = 30;
			sine[1768] = 30;
			sine[1769] = 31;
			sine[1770] = 31;
			sine[1771] = 31;
			sine[1772] = 31;
			sine[1773] = 32;
			sine[1774] = 32;
			sine[1775] = 32;
			sine[1776] = 32;
			sine[1777] = 33;
			sine[1778] = 33;
			sine[1779] = 33;
			sine[1780] = 33;
			sine[1781] = 34;
			sine[1782] = 34;
			sine[1783] = 34;
			sine[1784] = 35;
			sine[1785] = 35;
			sine[1786] = 35;
			sine[1787] = 35;
			sine[1788] = 36;
			sine[1789] = 36;
			sine[1790] = 36;
			sine[1791] = 36;
			sine[1792] = 37;
			sine[1793] = 37;
			sine[1794] = 37;
			sine[1795] = 38;
			sine[1796] = 38;
			sine[1797] = 38;
			sine[1798] = 38;
			sine[1799] = 39;
			sine[1800] = 39;
			sine[1801] = 39;
			sine[1802] = 39;
			sine[1803] = 40;
			sine[1804] = 40;
			sine[1805] = 40;
			sine[1806] = 41;
			sine[1807] = 41;
			sine[1808] = 41;
			sine[1809] = 42;
			sine[1810] = 42;
			sine[1811] = 42;
			sine[1812] = 42;
			sine[1813] = 43;
			sine[1814] = 43;
			sine[1815] = 43;
			sine[1816] = 44;
			sine[1817] = 44;
			sine[1818] = 44;
			sine[1819] = 44;
			sine[1820] = 45;
			sine[1821] = 45;
			sine[1822] = 45;
			sine[1823] = 46;
			sine[1824] = 46;
			sine[1825] = 46;
			sine[1826] = 47;
			sine[1827] = 47;
			sine[1828] = 47;
			sine[1829] = 47;
			sine[1830] = 48;
			sine[1831] = 48;
			sine[1832] = 48;
			sine[1833] = 49;
			sine[1834] = 49;
			sine[1835] = 49;
			sine[1836] = 50;
			sine[1837] = 50;
			sine[1838] = 50;
			sine[1839] = 51;
			sine[1840] = 51;
			sine[1841] = 51;
			sine[1842] = 51;
			sine[1843] = 52;
			sine[1844] = 52;
			sine[1845] = 52;
			sine[1846] = 53;
			sine[1847] = 53;
			sine[1848] = 53;
			sine[1849] = 54;
			sine[1850] = 54;
			sine[1851] = 54;
			sine[1852] = 55;
			sine[1853] = 55;
			sine[1854] = 55;
			sine[1855] = 56;
			sine[1856] = 56;
			sine[1857] = 56;
			sine[1858] = 57;
			sine[1859] = 57;
			sine[1860] = 57;
			sine[1861] = 58;
			sine[1862] = 58;
			sine[1863] = 58;
			sine[1864] = 59;
			sine[1865] = 59;
			sine[1866] = 59;
			sine[1867] = 60;
			sine[1868] = 60;
			sine[1869] = 60;
			sine[1870] = 61;
			sine[1871] = 61;
			sine[1872] = 61;
			sine[1873] = 62;
			sine[1874] = 62;
			sine[1875] = 62;
			sine[1876] = 63;
			sine[1877] = 63;
			sine[1878] = 63;
			sine[1879] = 64;
			sine[1880] = 64;
			sine[1881] = 64;
			sine[1882] = 65;
			sine[1883] = 65;
			sine[1884] = 65;
			sine[1885] = 66;
			sine[1886] = 66;
			sine[1887] = 66;
			sine[1888] = 67;
			sine[1889] = 67;
			sine[1890] = 67;
			sine[1891] = 68;
			sine[1892] = 68;
			sine[1893] = 68;
			sine[1894] = 69;
			sine[1895] = 69;
			sine[1896] = 69;
			sine[1897] = 70;
			sine[1898] = 70;
			sine[1899] = 70;
			sine[1900] = 71;
			sine[1901] = 71;
			sine[1902] = 71;
			sine[1903] = 72;
			sine[1904] = 72;
			sine[1905] = 73;
			sine[1906] = 73;
			sine[1907] = 73;
			sine[1908] = 74;
			sine[1909] = 74;
			sine[1910] = 74;
			sine[1911] = 75;
			sine[1912] = 75;
			sine[1913] = 75;
			sine[1914] = 76;
			sine[1915] = 76;
			sine[1916] = 76;
			sine[1917] = 77;
			sine[1918] = 77;
			sine[1919] = 78;
			sine[1920] = 78;
			sine[1921] = 78;
			sine[1922] = 79;
			sine[1923] = 79;
			sine[1924] = 79;
			sine[1925] = 80;
			sine[1926] = 80;
			sine[1927] = 80;
			sine[1928] = 81;
			sine[1929] = 81;
			sine[1930] = 82;
			sine[1931] = 82;
			sine[1932] = 82;
			sine[1933] = 83;
			sine[1934] = 83;
			sine[1935] = 83;
			sine[1936] = 84;
			sine[1937] = 84;
			sine[1938] = 84;
			sine[1939] = 85;
			sine[1940] = 85;
			sine[1941] = 86;
			sine[1942] = 86;
			sine[1943] = 86;
			sine[1944] = 87;
			sine[1945] = 87;
			sine[1946] = 87;
			sine[1947] = 88;
			sine[1948] = 88;
			sine[1949] = 89;
			sine[1950] = 89;
			sine[1951] = 89;
			sine[1952] = 90;
			sine[1953] = 90;
			sine[1954] = 90;
			sine[1955] = 91;
			sine[1956] = 91;
			sine[1957] = 92;
			sine[1958] = 92;
			sine[1959] = 92;
			sine[1960] = 93;
			sine[1961] = 93;
			sine[1962] = 93;
			sine[1963] = 94;
			sine[1964] = 94;
			sine[1965] = 95;
			sine[1966] = 95;
			sine[1967] = 95;
			sine[1968] = 96;
			sine[1969] = 96;
			sine[1970] = 96;
			sine[1971] = 97;
			sine[1972] = 97;
			sine[1973] = 98;
			sine[1974] = 98;
			sine[1975] = 98;
			sine[1976] = 99;
			sine[1977] = 99;
			sine[1978] = 99;
			sine[1979] = 100;
			sine[1980] = 100;
			sine[1981] = 101;
			sine[1982] = 101;
			sine[1983] = 101;
			sine[1984] = 102;
			sine[1985] = 102;
			sine[1986] = 102;
			sine[1987] = 103;
			sine[1988] = 103;
			sine[1989] = 104;
			sine[1990] = 104;
			sine[1991] = 104;
			sine[1992] = 105;
			sine[1993] = 105;
			sine[1994] = 106;
			sine[1995] = 106;
			sine[1996] = 106;
			sine[1997] = 107;
			sine[1998] = 107;
			sine[1999] = 107;
			sine[2000] = 108;
			sine[2001] = 108;
			sine[2002] = 109;
			sine[2003] = 109;
			sine[2004] = 109;
			sine[2005] = 110;
			sine[2006] = 110;
			sine[2007] = 111;
			sine[2008] = 111;
			sine[2009] = 111;
			sine[2010] = 112;
			sine[2011] = 112;
			sine[2012] = 113;
			sine[2013] = 113;
			sine[2014] = 113;
			sine[2015] = 114;
			sine[2016] = 114;
			sine[2017] = 114;
			sine[2018] = 115;
			sine[2019] = 115;
			sine[2020] = 116;
			sine[2021] = 116;
			sine[2022] = 116;
			sine[2023] = 117;
			sine[2024] = 117;
			sine[2025] = 118;
			sine[2026] = 118;
			sine[2027] = 118;
			sine[2028] = 119;
			sine[2029] = 119;
			sine[2030] = 119;
			sine[2031] = 120;
			sine[2032] = 120;
			sine[2033] = 121;
			sine[2034] = 121;
			sine[2035] = 121;
			sine[2036] = 122;
			sine[2037] = 122;
			sine[2038] = 123;
			sine[2039] = 123;
			sine[2040] = 123;
			sine[2041] = 124;
			sine[2042] = 124;
			sine[2043] = 125;
			sine[2044] = 125;
			sine[2045] = 125;
			sine[2046] = 126;
			sine[2047] = 126;
		end
endmodule
