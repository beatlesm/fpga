module input_signal_cos(radio_clk, codeword0, codeword1,codeword2,codeword3, codeword4, codeword5, codeword6, codeword7,codeword8, codeword9, codeword10, codeword11, codeword12, codeword13, codeword14, codeword15, codeword16, codeword17, codeword18, codeword19, codeword20, codeword21, codeword22, codeword23, codeword24, codeword25, codeword26, codeword27, codeword28, codeword29, codeword30, codeword31, codeword32, codeword33, codeword34, codeword35, codeword36, codeword37, codeword38, codeword39, codeword40, codeword41, codeword42, codeword43, codeword44, codeword45, codeword46, codeword47, codeword48, codeword49, get_tx);
//
	input radio_clk;
	input [31:0] codeword0, codeword1, codeword2, codeword3, codeword4,codeword5, codeword6,codeword7, codeword8, codeword9, codeword10, codeword11, codeword12, codeword13, codeword14, codeword15, codeword16, codeword17, codeword18, codeword19, codeword20, codeword21, codeword22, codeword23, codeword24, codeword25, codeword26, codeword27, codeword28, codeword29, codeword30, codeword31, codeword32, codeword33, codeword34, codeword35, codeword36, codeword37, codeword38, codeword39, codeword40, codeword41, codeword42, codeword43, codeword44, codeword45, codeword46, codeword47, codeword48, codeword49;

   output [31:0] get_tx;

	reg [15:0] phase_acc0, phase_acc1, phase_acc2, phase_acc3, phase_acc4, phase_acc5, phase_acc6, phase_acc7, phase_acc8, phase_acc9, phase_acc10, phase_acc11, phase_acc12, phase_acc13, phase_acc14, phase_acc15, phase_acc16, phase_acc17, phase_acc18, phase_acc19, phase_acc20, phase_acc21, phase_acc22, phase_acc23, phase_acc24, phase_acc25, phase_acc26, phase_acc27, phase_acc28, phase_acc29, phase_acc30, phase_acc31, phase_acc32, phase_acc33, phase_acc34, phase_acc35, phase_acc36, phase_acc37, phase_acc38, phase_acc39, phase_acc40, phase_acc41, phase_acc42, phase_acc43, phase_acc44, phase_acc45, phase_acc46, phase_acc47, phase_acc48, phase_acc49;

   reg [31:0] tx_out;

   reg [15:0] freq0, freq1, freq2, freq3, freq4, freq5, freq6, freq7, freq8, freq9, freq10, freq11, freq12, freq13, freq14, freq15, freq16, freq17, freq18, freq19, freq20, freq21, freq22, freq23, freq24, freq25, freq26, freq27, freq28, freq29, freq30, freq31, freq32, freq33, freq34, freq35, freq36, freq37, freq38, freq39, freq40, freq41, freq42, freq43, freq44, freq45, freq46, freq47, freq48, freq49;
	reg [7:0] amp0, amp1, amp2, amp3, amp4, amp5, amp6, amp7, amp8, amp9, amp10, amp11, amp12, amp13, amp14, amp15, amp16, amp17, amp18, amp19, amp20, amp21, amp22, amp23, amp24, amp25, amp26, amp27, amp28, amp29, amp30, amp31, amp32, amp33, amp34, amp35, amp36, amp37, amp38, amp39, amp40, amp41, amp42, amp43, amp44, amp45, amp46, amp47, amp48, amp49;
   reg [10:0] ph0, ph1, ph2, ph3, ph4, ph5, ph6, ph7, ph8, ph9, ph10, ph11, ph12, ph13, ph14, ph15, ph16, ph17, ph18, ph19, ph20, ph21, ph22, ph23, ph24, ph25, ph26, ph27, ph28, ph29, ph30, ph31, ph32, ph33, ph34, ph35, ph36, ph37, ph38, ph39, ph40, ph41, ph42, ph43, ph44, ph45, ph46, ph47, ph48, ph49;
   reg [7:0] tmp;

	reg [25:0] amp_times_sin; // 26 bits: 8 bits for amplitude, 10 bits for sine wave, 6 bits for 50 frequencies, and two bits for coercion
	reg [15:0] neg_amp_times_sin;
	
    always @(posedge radio_clk) begin

			freq0 = codeword0[15:0];
			amp0 = codeword0[23:16];
			tmp=codeword0[31:24];
			ph0 = tmp << 3;

			freq1 = codeword1[15:0];
			amp1 = codeword1[23:16];
			tmp=codeword1[31:24];
			ph1 = tmp << 3;

			freq2 = codeword2[15:0];
			amp2 = codeword2[23:16];
			tmp=codeword2[31:24];
			ph2 = tmp << 3;

			freq3 = codeword3[15:0];
			amp3 = codeword3[23:16];
			tmp=codeword3[31:24];
			ph3 = tmp << 3;

			freq4 = codeword4[15:0];
			amp4 = codeword4[23:16];
			tmp=codeword4[31:24];
			ph4 = tmp << 3;

			freq5 = codeword5[15:0];
			amp5 = codeword5[23:16];
			tmp=codeword5[31:24];
			ph5 = tmp << 3;

			freq6 = codeword6[15:0];
			amp6 = codeword6[23:16];
			tmp=codeword6[31:24];
			ph6 = tmp << 3;

			freq7 = codeword7[15:0];
			amp7 = codeword7[23:16];
			tmp=codeword7[31:24];
			ph7 = tmp << 3;

			freq8 = codeword8[15:0];
			amp8 = codeword8[23:16];
			tmp=codeword8[31:24];
			ph8 = tmp << 3;

			freq9 = codeword9[15:0];
			amp9 = codeword9[23:16];
			tmp=codeword9[31:24];
			ph9 = tmp << 3;

			freq10 = codeword10[15:0];
			amp10 = codeword10[23:16];
			tmp=codeword10[31:24];
			ph10 = tmp << 3;

			freq11 = codeword11[15:0];
			amp11 = codeword11[23:16];
			tmp=codeword11[31:24];
			ph11 = tmp << 3;

			freq12 = codeword12[15:0];
			amp12 = codeword12[23:16];
			tmp=codeword12[31:24];
			ph12 = tmp << 3;

			freq13 = codeword13[15:0];
			amp13 = codeword13[23:16];
			tmp=codeword13[31:24];
			ph13 = tmp << 3;

			freq14 = codeword14[15:0];
			amp14 = codeword14[23:16];
			tmp=codeword14[31:24];
			ph14 = tmp << 3;

			freq15 = codeword15[15:0];
			amp15 = codeword15[23:16];
			tmp=codeword15[31:24];
			ph15 = tmp << 3;

			freq16 = codeword16[15:0];
			amp16 = codeword16[23:16];
			tmp=codeword16[31:24];
			ph16 = tmp << 3;

			freq17 = codeword17[15:0];
			amp17 = codeword17[23:16];
			tmp=codeword17[31:24];
			ph17 = tmp << 3;

			freq18 = codeword18[15:0];
			amp18 = codeword18[23:16];
			tmp=codeword18[31:24];
			ph18 = tmp << 3;

			freq19 = codeword19[15:0];
			amp19 = codeword19[23:16];
			tmp=codeword19[31:24];
			ph19 = tmp << 3;

			freq20 = codeword20[15:0];
			amp20 = codeword20[23:16];
			tmp = codeword20[31:24];
			ph20 = tmp << 3;

			freq21 = codeword21[15:0];
			amp21 = codeword21[23:16];
			tmp = codeword21[31:24];
			ph21 = tmp << 3;

			freq22 = codeword22[15:0];
			amp22 = codeword22[23:16];
			tmp = codeword22[31:24];
			ph22 = tmp << 3;

			freq23 = codeword23[15:0];
			amp23 = codeword23[23:16];
			tmp = codeword23[31:24];
			ph23 = tmp << 3;

			freq24 = codeword24[15:0];
			amp24 = codeword24[23:16];
			tmp = codeword24[31:24];
			ph24 = tmp << 3;

			freq25 = codeword25[15:0];
			amp25 = codeword25[23:16];
			tmp = codeword25[31:24];
			ph25 = tmp << 3;

			freq26 = codeword26[15:0];
			amp26 = codeword26[23:16];
			tmp = codeword26[31:24];
			ph26 = tmp << 3;

			freq27 = codeword27[15:0];
			amp27 = codeword27[23:16];
			tmp = codeword27[31:24];
			ph27 = tmp << 3;

			freq28 = codeword28[15:0];
			amp28 = codeword28[23:16];
			tmp = codeword28[31:24];
			ph28 = tmp << 3;

			freq29 = codeword29[15:0];
			amp29 = codeword29[23:16];
			tmp = codeword29[31:24];
			ph29 = tmp << 3;

			freq30 = codeword30[15:0];
			amp30 = codeword30[23:16];
			tmp = codeword30[31:24];
			ph30 = tmp << 3;

			freq31 = codeword31[15:0];
			amp31 = codeword31[23:16];
			tmp = codeword31[31:24];
			ph31 = tmp << 3;

			freq32 = codeword32[15:0];
			amp32 = codeword32[23:16];
			tmp = codeword32[31:24];
			ph32 = tmp << 3;

			freq33 = codeword33[15:0];
			amp33 = codeword33[23:16];
			tmp = codeword33[31:24];
			ph33 = tmp << 3;

			freq34 = codeword34[15:0];
			amp34 = codeword34[23:16];
			tmp = codeword34[31:24];
			ph34 = tmp << 3;

			freq35 = codeword35[15:0];
			amp35 = codeword35[23:16];
			tmp = codeword35[31:24];
			ph35 = tmp << 3;

			freq36 = codeword36[15:0];
			amp36 = codeword36[23:16];
			tmp = codeword36[31:24];
			ph36 = tmp << 3;

			freq37 = codeword37[15:0];
			amp37 = codeword37[23:16];
			tmp = codeword37[31:24];
			ph37 = tmp << 3;

			freq38 = codeword38[15:0];
			amp38 = codeword38[23:16];
			tmp = codeword38[31:24];
			ph38 = tmp << 3;

			freq39 = codeword39[15:0];
			amp39 = codeword39[23:16];
			tmp = codeword39[31:24];
			ph39 = tmp << 3;

			freq40 = codeword40[15:0];
			amp40 = codeword40[23:16];
			tmp = codeword40[31:24];
			ph40 = tmp << 3;

			freq41 = codeword41[15:0];
			amp41 = codeword41[23:16];
			tmp = codeword41[31:24];
			ph41 = tmp << 3;

			freq42 = codeword42[15:0];
			amp42 = codeword42[23:16];
			tmp = codeword42[31:24];
			ph42 = tmp << 3;

			freq43 = codeword43[15:0];
			amp43 = codeword43[23:16];
			tmp = codeword43[31:24];
			ph43 = tmp << 3;

			freq44 = codeword44[15:0];
			amp44 = codeword44[23:16];
			tmp = codeword44[31:24];
			ph44 = tmp << 3;

			freq45 = codeword45[15:0];
			amp45 = codeword45[23:16];
			tmp = codeword45[31:24];
			ph45 = tmp << 3;

			freq46 = codeword46[15:0];
			amp46 = codeword46[23:16];
			tmp = codeword46[31:24];
			ph46 = tmp << 3;

			freq47 = codeword47[15:0];
			amp47 = codeword47[23:16];
			tmp = codeword47[31:24];
			ph47 = tmp << 3;

			freq48 = codeword48[15:0];
			amp48 = codeword48[23:16];
			tmp = codeword48[31:24];
			ph48 = tmp << 3;

			freq49 = codeword49[15:0];
			amp49 = codeword49[23:16];
			tmp = codeword49[31:24];
			ph49 = tmp << 3;
			phase_acc0 = phase_acc0 + freq0;
			phase_acc1 = phase_acc1 + freq1;
			phase_acc2 = phase_acc2 + freq2;
			phase_acc3 = phase_acc3 + freq3;
			phase_acc4 = phase_acc4 + freq4;
			phase_acc5 = phase_acc5 + freq5;
			phase_acc6 = phase_acc6 + freq6;
			phase_acc7 = phase_acc7 + freq7;
			phase_acc8 = phase_acc8 + freq8;
			phase_acc9 = phase_acc9 + freq9;
			phase_acc10 = phase_acc10 + freq10;
			phase_acc11 = phase_acc11 + freq11;
			phase_acc12 = phase_acc12 + freq12;
			phase_acc13 = phase_acc13 + freq13;
			phase_acc14 = phase_acc14 + freq14;
			phase_acc15 = phase_acc15 + freq15;
			phase_acc16 = phase_acc16 + freq16;
			phase_acc17 = phase_acc17 + freq17;
			phase_acc18 = phase_acc18 + freq18;
			phase_acc19 = phase_acc19 + freq19;
			phase_acc20 = phase_acc20 + freq20;
			phase_acc21 = phase_acc21 + freq21;
			phase_acc22 = phase_acc22 + freq22;
			phase_acc23 = phase_acc23 + freq23;
			phase_acc24 = phase_acc24 + freq24;
			phase_acc25 = phase_acc25 + freq25;
			phase_acc26 = phase_acc26 + freq26;
			phase_acc27 = phase_acc27 + freq27;
			phase_acc28 = phase_acc28 + freq28;
			phase_acc29 = phase_acc29 + freq29;
			phase_acc30 = phase_acc30 + freq30;
			phase_acc31 = phase_acc31 + freq31;
			phase_acc32 = phase_acc32 + freq32;
			phase_acc33 = phase_acc33 + freq33;
			phase_acc34 = phase_acc34 + freq34;
			phase_acc35 = phase_acc35 + freq35;
			phase_acc36 = phase_acc36 + freq36;
			phase_acc37 = phase_acc37 + freq37;
			phase_acc38 = phase_acc38 + freq38;
			phase_acc39 = phase_acc39 + freq39;
			phase_acc40 = phase_acc40 + freq40;
			phase_acc41 = phase_acc41 + freq41;
			phase_acc42 = phase_acc42 + freq42;
			phase_acc43 = phase_acc43 + freq43;
			phase_acc44 = phase_acc44 + freq44;
			phase_acc45 = phase_acc45 + freq45;
			phase_acc46 = phase_acc46 + freq46;
			phase_acc47 = phase_acc47 + freq47;
			phase_acc48 = phase_acc48 + freq48;
			phase_acc49 = phase_acc49 + freq49;
		amp_times_sin = amp0*cos[phase_acc0[15:5] + ph0] + amp1*cos[phase_acc1[15:5] + ph1] + amp2*cos[phase_acc2[15:5] + ph2] + amp3*cos[phase_acc3[15:5] + ph3] + amp4*cos[phase_acc4[15:5] + ph4] + amp5*cos[phase_acc5[15:5] + ph5] + amp6*cos[phase_acc6[15:5] + ph6] + amp7*cos[phase_acc7[15:5] + ph7] + amp8*cos[phase_acc8[15:5] + ph8] + amp9*cos[phase_acc9[15:5] + ph9] + amp10*cos[phase_acc10[15:5] + ph10] + amp11*cos[phase_acc11[15:5] + ph11] + amp12*cos[phase_acc12[15:5] + ph12] + amp13*cos[phase_acc13[15:5] + ph13] + amp14*cos[phase_acc14[15:5] + ph14] + amp15*cos[phase_acc15[15:5] + ph15] + amp16*cos[phase_acc16[15:5] + ph16] + amp17*cos[phase_acc17[15:5] + ph17] + amp18*cos[phase_acc18[15:5] + ph18] + amp19*cos[phase_acc19[15:5] + ph19];// + amp20*cos[phase_acc20[15:5] + ph20] + amp21*cos[phase_acc21[15:5] + ph21] + amp22*cos[phase_acc22[15:5] + ph22] + amp23*cos[phase_acc23[15:5] + ph23] + amp24*cos[phase_acc24[15:5] + ph24] + amp25*cos[phase_acc25[15:5] + ph25] + amp26*cos[phase_acc26[15:5] + ph26] + amp27*cos[phase_acc27[15:5] + ph27] + amp28*cos[phase_acc28[15:5] + ph28] + amp29*cos[phase_acc29[15:5] + ph29] + amp30*cos[phase_acc30[15:5] + ph30] + amp31*cos[phase_acc31[15:5] + ph31] + amp32*cos[phase_acc32[15:5] + ph32] + amp33*cos[phase_acc33[15:5] + ph33] + amp34*cos[phase_acc34[15:5] + ph34] + amp35*cos[phase_acc35[15:5] + ph35] + amp36*cos[phase_acc36[15:5] + ph36] + amp37*cos[phase_acc37[15:5] + ph37] + amp38*cos[phase_acc38[15:5] + ph38] + amp39*cos[phase_acc39[15:5] + ph39] + amp40*cos[phase_acc40[15:5] + ph40] + amp41*cos[phase_acc41[15:5] + ph41] + amp42*cos[phase_acc42[15:5] + ph42] + amp43*cos[phase_acc43[15:5] + ph43] + amp44*cos[phase_acc44[15:5] + ph44] + amp45*cos[phase_acc45[15:5] + ph45] + amp46*cos[phase_acc46[15:5] + ph46] + amp47*cos[phase_acc47[15:5] + ph47] + amp48*cos[phase_acc48[15:5] + ph48] + amp49*cos[phase_acc49[15:5] + ph49]; 

			tx_out[15:0] = amp_times_sin[23:8];
			begin
				if (amp_times_sin[25] == 1 || amp_times_sin[24] == 1) 
					tx_out[15:0] = 16'b1111111111111111; // Coercion line. 
			end
		  tx_out[31:16] = amp_times_sin[23:8];//16'b0000000000000000;
//        tx_out[31:16] = 16'b0000000000000000;
		  // Trying IQ channel thing
		//  tx_out[31:16] =  amp_times_sin[23:8];
		//   	tx[31:16] <= (run_tx) ? get_tx[31:16] : tx_idle[31:16]; // I channel

    end
   assign get_tx = tx_out;


// SINE LOOKUP TABLE
    reg [9:0] cos [0:2047];
    initial
        begin
				cos[0] = 682;
				cos[1] = 682;
				cos[2] = 682;
				cos[3] = 682;
				cos[4] = 682;
				cos[5] = 682;
				cos[6] = 682;
				cos[7] = 682;
				cos[8] = 682;
				cos[9] = 682;
				cos[10] = 682;
				cos[11] = 682;
				cos[12] = 682;
				cos[13] = 682;
				cos[14] = 682;
				cos[15] = 682;
				cos[16] = 682;
				cos[17] = 682;
				cos[18] = 682;
				cos[19] = 682;
				cos[20] = 682;
				cos[21] = 681;
				cos[22] = 681;
				cos[23] = 681;
				cos[24] = 681;
				cos[25] = 681;
				cos[26] = 681;
				cos[27] = 681;
				cos[28] = 681;
				cos[29] = 681;
				cos[30] = 681;
				cos[31] = 681;
				cos[32] = 681;
				cos[33] = 680;
				cos[34] = 680;
				cos[35] = 680;
				cos[36] = 680;
				cos[37] = 680;
				cos[38] = 680;
				cos[39] = 680;
				cos[40] = 680;
				cos[41] = 679;
				cos[42] = 679;
				cos[43] = 679;
				cos[44] = 679;
				cos[45] = 679;
				cos[46] = 679;
				cos[47] = 679;
				cos[48] = 678;
				cos[49] = 678;
				cos[50] = 678;
				cos[51] = 678;
				cos[52] = 678;
				cos[53] = 678;
				cos[54] = 677;
				cos[55] = 677;
				cos[56] = 677;
				cos[57] = 677;
				cos[58] = 677;
				cos[59] = 677;
				cos[60] = 676;
				cos[61] = 676;
				cos[62] = 676;
				cos[63] = 676;
				cos[64] = 676;
				cos[65] = 675;
				cos[66] = 675;
				cos[67] = 675;
				cos[68] = 675;
				cos[69] = 675;
				cos[70] = 674;
				cos[71] = 674;
				cos[72] = 674;
				cos[73] = 674;
				cos[74] = 673;
				cos[75] = 673;
				cos[76] = 673;
				cos[77] = 673;
				cos[78] = 672;
				cos[79] = 672;
				cos[80] = 672;
				cos[81] = 672;
				cos[82] = 671;
				cos[83] = 671;
				cos[84] = 671;
				cos[85] = 671;
				cos[86] = 670;
				cos[87] = 670;
				cos[88] = 670;
				cos[89] = 670;
				cos[90] = 669;
				cos[91] = 669;
				cos[92] = 669;
				cos[93] = 668;
				cos[94] = 668;
				cos[95] = 668;
				cos[96] = 667;
				cos[97] = 667;
				cos[98] = 667;
				cos[99] = 667;
				cos[100] = 666;
				cos[101] = 666;
				cos[102] = 666;
				cos[103] = 665;
				cos[104] = 665;
				cos[105] = 665;
				cos[106] = 664;
				cos[107] = 664;
				cos[108] = 664;
				cos[109] = 663;
				cos[110] = 663;
				cos[111] = 663;
				cos[112] = 662;
				cos[113] = 662;
				cos[114] = 662;
				cos[115] = 661;
				cos[116] = 661;
				cos[117] = 660;
				cos[118] = 660;
				cos[119] = 660;
				cos[120] = 659;
				cos[121] = 659;
				cos[122] = 659;
				cos[123] = 658;
				cos[124] = 658;
				cos[125] = 657;
				cos[126] = 657;
				cos[127] = 657;
				cos[128] = 656;
				cos[129] = 656;
				cos[130] = 655;
				cos[131] = 655;
				cos[132] = 655;
				cos[133] = 654;
				cos[134] = 654;
				cos[135] = 653;
				cos[136] = 653;
				cos[137] = 652;
				cos[138] = 652;
				cos[139] = 652;
				cos[140] = 651;
				cos[141] = 651;
				cos[142] = 650;
				cos[143] = 650;
				cos[144] = 649;
				cos[145] = 649;
				cos[146] = 648;
				cos[147] = 648;
				cos[148] = 648;
				cos[149] = 647;
				cos[150] = 647;
				cos[151] = 646;
				cos[152] = 646;
				cos[153] = 645;
				cos[154] = 645;
				cos[155] = 644;
				cos[156] = 644;
				cos[157] = 643;
				cos[158] = 643;
				cos[159] = 642;
				cos[160] = 642;
				cos[161] = 641;
				cos[162] = 641;
				cos[163] = 640;
				cos[164] = 640;
				cos[165] = 639;
				cos[166] = 639;
				cos[167] = 638;
				cos[168] = 638;
				cos[169] = 637;
				cos[170] = 637;
				cos[171] = 636;
				cos[172] = 636;
				cos[173] = 635;
				cos[174] = 635;
				cos[175] = 634;
				cos[176] = 634;
				cos[177] = 633;
				cos[178] = 633;
				cos[179] = 632;
				cos[180] = 631;
				cos[181] = 631;
				cos[182] = 630;
				cos[183] = 630;
				cos[184] = 629;
				cos[185] = 629;
				cos[186] = 628;
				cos[187] = 628;
				cos[188] = 627;
				cos[189] = 626;
				cos[190] = 626;
				cos[191] = 625;
				cos[192] = 625;
				cos[193] = 624;
				cos[194] = 623;
				cos[195] = 623;
				cos[196] = 622;
				cos[197] = 622;
				cos[198] = 621;
				cos[199] = 621;
				cos[200] = 620;
				cos[201] = 619;
				cos[202] = 619;
				cos[203] = 618;
				cos[204] = 617;
				cos[205] = 617;
				cos[206] = 616;
				cos[207] = 616;
				cos[208] = 615;
				cos[209] = 614;
				cos[210] = 614;
				cos[211] = 613;
				cos[212] = 612;
				cos[213] = 612;
				cos[214] = 611;
				cos[215] = 611;
				cos[216] = 610;
				cos[217] = 609;
				cos[218] = 609;
				cos[219] = 608;
				cos[220] = 607;
				cos[221] = 607;
				cos[222] = 606;
				cos[223] = 605;
				cos[224] = 605;
				cos[225] = 604;
				cos[226] = 603;
				cos[227] = 603;
				cos[228] = 602;
				cos[229] = 601;
				cos[230] = 601;
				cos[231] = 600;
				cos[232] = 599;
				cos[233] = 599;
				cos[234] = 598;
				cos[235] = 597;
				cos[236] = 597;
				cos[237] = 596;
				cos[238] = 595;
				cos[239] = 594;
				cos[240] = 594;
				cos[241] = 593;
				cos[242] = 592;
				cos[243] = 592;
				cos[244] = 591;
				cos[245] = 590;
				cos[246] = 589;
				cos[247] = 589;
				cos[248] = 588;
				cos[249] = 587;
				cos[250] = 587;
				cos[251] = 586;
				cos[252] = 585;
				cos[253] = 584;
				cos[254] = 584;
				cos[255] = 583;
				cos[256] = 582;
				cos[257] = 581;
				cos[258] = 581;
				cos[259] = 580;
				cos[260] = 579;
				cos[261] = 578;
				cos[262] = 578;
				cos[263] = 577;
				cos[264] = 576;
				cos[265] = 575;
				cos[266] = 575;
				cos[267] = 574;
				cos[268] = 573;
				cos[269] = 572;
				cos[270] = 572;
				cos[271] = 571;
				cos[272] = 570;
				cos[273] = 569;
				cos[274] = 569;
				cos[275] = 568;
				cos[276] = 567;
				cos[277] = 566;
				cos[278] = 565;
				cos[279] = 565;
				cos[280] = 564;
				cos[281] = 563;
				cos[282] = 562;
				cos[283] = 561;
				cos[284] = 561;
				cos[285] = 560;
				cos[286] = 559;
				cos[287] = 558;
				cos[288] = 557;
				cos[289] = 557;
				cos[290] = 556;
				cos[291] = 555;
				cos[292] = 554;
				cos[293] = 553;
				cos[294] = 552;
				cos[295] = 552;
				cos[296] = 551;
				cos[297] = 550;
				cos[298] = 549;
				cos[299] = 548;
				cos[300] = 548;
				cos[301] = 547;
				cos[302] = 546;
				cos[303] = 545;
				cos[304] = 544;
				cos[305] = 543;
				cos[306] = 542;
				cos[307] = 542;
				cos[308] = 541;
				cos[309] = 540;
				cos[310] = 539;
				cos[311] = 538;
				cos[312] = 537;
				cos[313] = 537;
				cos[314] = 536;
				cos[315] = 535;
				cos[316] = 534;
				cos[317] = 533;
				cos[318] = 532;
				cos[319] = 531;
				cos[320] = 530;
				cos[321] = 530;
				cos[322] = 529;
				cos[323] = 528;
				cos[324] = 527;
				cos[325] = 526;
				cos[326] = 525;
				cos[327] = 524;
				cos[328] = 523;
				cos[329] = 523;
				cos[330] = 522;
				cos[331] = 521;
				cos[332] = 520;
				cos[333] = 519;
				cos[334] = 518;
				cos[335] = 517;
				cos[336] = 516;
				cos[337] = 515;
				cos[338] = 515;
				cos[339] = 514;
				cos[340] = 513;
				cos[341] = 512;
				cos[342] = 511;
				cos[343] = 510;
				cos[344] = 509;
				cos[345] = 508;
				cos[346] = 507;
				cos[347] = 506;
				cos[348] = 505;
				cos[349] = 505;
				cos[350] = 504;
				cos[351] = 503;
				cos[352] = 502;
				cos[353] = 501;
				cos[354] = 500;
				cos[355] = 499;
				cos[356] = 498;
				cos[357] = 497;
				cos[358] = 496;
				cos[359] = 495;
				cos[360] = 494;
				cos[361] = 493;
				cos[362] = 492;
				cos[363] = 491;
				cos[364] = 491;
				cos[365] = 490;
				cos[366] = 489;
				cos[367] = 488;
				cos[368] = 487;
				cos[369] = 486;
				cos[370] = 485;
				cos[371] = 484;
				cos[372] = 483;
				cos[373] = 482;
				cos[374] = 481;
				cos[375] = 480;
				cos[376] = 479;
				cos[377] = 478;
				cos[378] = 477;
				cos[379] = 476;
				cos[380] = 475;
				cos[381] = 474;
				cos[382] = 473;
				cos[383] = 472;
				cos[384] = 471;
				cos[385] = 470;
				cos[386] = 470;
				cos[387] = 469;
				cos[388] = 468;
				cos[389] = 467;
				cos[390] = 466;
				cos[391] = 465;
				cos[392] = 464;
				cos[393] = 463;
				cos[394] = 462;
				cos[395] = 461;
				cos[396] = 460;
				cos[397] = 459;
				cos[398] = 458;
				cos[399] = 457;
				cos[400] = 456;
				cos[401] = 455;
				cos[402] = 454;
				cos[403] = 453;
				cos[404] = 452;
				cos[405] = 451;
				cos[406] = 450;
				cos[407] = 449;
				cos[408] = 448;
				cos[409] = 447;
				cos[410] = 446;
				cos[411] = 445;
				cos[412] = 444;
				cos[413] = 443;
				cos[414] = 442;
				cos[415] = 441;
				cos[416] = 440;
				cos[417] = 439;
				cos[418] = 438;
				cos[419] = 437;
				cos[420] = 436;
				cos[421] = 435;
				cos[422] = 434;
				cos[423] = 433;
				cos[424] = 432;
				cos[425] = 431;
				cos[426] = 430;
				cos[427] = 429;
				cos[428] = 428;
				cos[429] = 427;
				cos[430] = 426;
				cos[431] = 425;
				cos[432] = 424;
				cos[433] = 423;
				cos[434] = 422;
				cos[435] = 421;
				cos[436] = 420;
				cos[437] = 419;
				cos[438] = 418;
				cos[439] = 417;
				cos[440] = 416;
				cos[441] = 415;
				cos[442] = 414;
				cos[443] = 413;
				cos[444] = 412;
				cos[445] = 411;
				cos[446] = 409;
				cos[447] = 408;
				cos[448] = 407;
				cos[449] = 406;
				cos[450] = 405;
				cos[451] = 404;
				cos[452] = 403;
				cos[453] = 402;
				cos[454] = 401;
				cos[455] = 400;
				cos[456] = 399;
				cos[457] = 398;
				cos[458] = 397;
				cos[459] = 396;
				cos[460] = 395;
				cos[461] = 394;
				cos[462] = 393;
				cos[463] = 392;
				cos[464] = 391;
				cos[465] = 390;
				cos[466] = 389;
				cos[467] = 388;
				cos[468] = 387;
				cos[469] = 386;
				cos[470] = 385;
				cos[471] = 384;
				cos[472] = 383;
				cos[473] = 382;
				cos[474] = 381;
				cos[475] = 379;
				cos[476] = 378;
				cos[477] = 377;
				cos[478] = 376;
				cos[479] = 375;
				cos[480] = 374;
				cos[481] = 373;
				cos[482] = 372;
				cos[483] = 371;
				cos[484] = 370;
				cos[485] = 369;
				cos[486] = 368;
				cos[487] = 367;
				cos[488] = 366;
				cos[489] = 365;
				cos[490] = 364;
				cos[491] = 363;
				cos[492] = 362;
				cos[493] = 361;
				cos[494] = 360;
				cos[495] = 359;
				cos[496] = 358;
				cos[497] = 357;
				cos[498] = 355;
				cos[499] = 354;
				cos[500] = 353;
				cos[501] = 352;
				cos[502] = 351;
				cos[503] = 350;
				cos[504] = 349;
				cos[505] = 348;
				cos[506] = 347;
				cos[507] = 346;
				cos[508] = 345;
				cos[509] = 344;
				cos[510] = 343;
				cos[511] = 342;
				cos[512] = 341;
				cos[513] = 340;
				cos[514] = 339;
				cos[515] = 338;
				cos[516] = 337;
				cos[517] = 336;
				cos[518] = 335;
				cos[519] = 334;
				cos[520] = 332;
				cos[521] = 331;
				cos[522] = 330;
				cos[523] = 329;
				cos[524] = 328;
				cos[525] = 327;
				cos[526] = 326;
				cos[527] = 325;
				cos[528] = 324;
				cos[529] = 323;
				cos[530] = 322;
				cos[531] = 321;
				cos[532] = 320;
				cos[533] = 319;
				cos[534] = 318;
				cos[535] = 317;
				cos[536] = 316;
				cos[537] = 315;
				cos[538] = 314;
				cos[539] = 313;
				cos[540] = 312;
				cos[541] = 311;
				cos[542] = 309;
				cos[543] = 308;
				cos[544] = 307;
				cos[545] = 306;
				cos[546] = 305;
				cos[547] = 304;
				cos[548] = 303;
				cos[549] = 302;
				cos[550] = 301;
				cos[551] = 300;
				cos[552] = 299;
				cos[553] = 298;
				cos[554] = 297;
				cos[555] = 296;
				cos[556] = 295;
				cos[557] = 294;
				cos[558] = 293;
				cos[559] = 292;
				cos[560] = 291;
				cos[561] = 290;
				cos[562] = 289;
				cos[563] = 288;
				cos[564] = 287;
				cos[565] = 286;
				cos[566] = 285;
				cos[567] = 284;
				cos[568] = 282;
				cos[569] = 281;
				cos[570] = 280;
				cos[571] = 279;
				cos[572] = 278;
				cos[573] = 277;
				cos[574] = 276;
				cos[575] = 275;
				cos[576] = 274;
				cos[577] = 273;
				cos[578] = 272;
				cos[579] = 271;
				cos[580] = 270;
				cos[581] = 269;
				cos[582] = 268;
				cos[583] = 267;
				cos[584] = 266;
				cos[585] = 265;
				cos[586] = 264;
				cos[587] = 263;
				cos[588] = 262;
				cos[589] = 261;
				cos[590] = 260;
				cos[591] = 259;
				cos[592] = 258;
				cos[593] = 257;
				cos[594] = 256;
				cos[595] = 255;
				cos[596] = 254;
				cos[597] = 253;
				cos[598] = 252;
				cos[599] = 251;
				cos[600] = 250;
				cos[601] = 249;
				cos[602] = 248;
				cos[603] = 247;
				cos[604] = 246;
				cos[605] = 245;
				cos[606] = 244;
				cos[607] = 243;
				cos[608] = 242;
				cos[609] = 241;
				cos[610] = 240;
				cos[611] = 239;
				cos[612] = 238;
				cos[613] = 237;
				cos[614] = 236;
				cos[615] = 235;
				cos[616] = 234;
				cos[617] = 233;
				cos[618] = 232;
				cos[619] = 231;
				cos[620] = 230;
				cos[621] = 229;
				cos[622] = 228;
				cos[623] = 227;
				cos[624] = 226;
				cos[625] = 225;
				cos[626] = 224;
				cos[627] = 223;
				cos[628] = 222;
				cos[629] = 221;
				cos[630] = 220;
				cos[631] = 219;
				cos[632] = 218;
				cos[633] = 217;
				cos[634] = 216;
				cos[635] = 215;
				cos[636] = 214;
				cos[637] = 213;
				cos[638] = 212;
				cos[639] = 211;
				cos[640] = 210;
				cos[641] = 209;
				cos[642] = 208;
				cos[643] = 207;
				cos[644] = 206;
				cos[645] = 205;
				cos[646] = 204;
				cos[647] = 203;
				cos[648] = 203;
				cos[649] = 202;
				cos[650] = 201;
				cos[651] = 200;
				cos[652] = 199;
				cos[653] = 198;
				cos[654] = 197;
				cos[655] = 196;
				cos[656] = 195;
				cos[657] = 194;
				cos[658] = 193;
				cos[659] = 192;
				cos[660] = 191;
				cos[661] = 190;
				cos[662] = 189;
				cos[663] = 188;
				cos[664] = 187;
				cos[665] = 186;
				cos[666] = 185;
				cos[667] = 185;
				cos[668] = 184;
				cos[669] = 183;
				cos[670] = 182;
				cos[671] = 181;
				cos[672] = 180;
				cos[673] = 179;
				cos[674] = 178;
				cos[675] = 177;
				cos[676] = 176;
				cos[677] = 175;
				cos[678] = 174;
				cos[679] = 174;
				cos[680] = 173;
				cos[681] = 172;
				cos[682] = 171;
				cos[683] = 170;
				cos[684] = 169;
				cos[685] = 168;
				cos[686] = 167;
				cos[687] = 166;
				cos[688] = 165;
				cos[689] = 164;
				cos[690] = 164;
				cos[691] = 163;
				cos[692] = 162;
				cos[693] = 161;
				cos[694] = 160;
				cos[695] = 159;
				cos[696] = 158;
				cos[697] = 157;
				cos[698] = 156;
				cos[699] = 156;
				cos[700] = 155;
				cos[701] = 154;
				cos[702] = 153;
				cos[703] = 152;
				cos[704] = 151;
				cos[705] = 150;
				cos[706] = 149;
				cos[707] = 149;
				cos[708] = 148;
				cos[709] = 147;
				cos[710] = 146;
				cos[711] = 145;
				cos[712] = 144;
				cos[713] = 143;
				cos[714] = 143;
				cos[715] = 142;
				cos[716] = 141;
				cos[717] = 140;
				cos[718] = 139;
				cos[719] = 138;
				cos[720] = 138;
				cos[721] = 137;
				cos[722] = 136;
				cos[723] = 135;
				cos[724] = 134;
				cos[725] = 133;
				cos[726] = 132;
				cos[727] = 132;
				cos[728] = 131;
				cos[729] = 130;
				cos[730] = 129;
				cos[731] = 128;
				cos[732] = 128;
				cos[733] = 127;
				cos[734] = 126;
				cos[735] = 125;
				cos[736] = 124;
				cos[737] = 123;
				cos[738] = 123;
				cos[739] = 122;
				cos[740] = 121;
				cos[741] = 120;
				cos[742] = 119;
				cos[743] = 119;
				cos[744] = 118;
				cos[745] = 117;
				cos[746] = 116;
				cos[747] = 116;
				cos[748] = 115;
				cos[749] = 114;
				cos[750] = 113;
				cos[751] = 112;
				cos[752] = 112;
				cos[753] = 111;
				cos[754] = 110;
				cos[755] = 109;
				cos[756] = 109;
				cos[757] = 108;
				cos[758] = 107;
				cos[759] = 106;
				cos[760] = 105;
				cos[761] = 105;
				cos[762] = 104;
				cos[763] = 103;
				cos[764] = 102;
				cos[765] = 102;
				cos[766] = 101;
				cos[767] = 100;
				cos[768] = 99;
				cos[769] = 99;
				cos[770] = 98;
				cos[771] = 97;
				cos[772] = 97;
				cos[773] = 96;
				cos[774] = 95;
				cos[775] = 94;
				cos[776] = 94;
				cos[777] = 93;
				cos[778] = 92;
				cos[779] = 91;
				cos[780] = 91;
				cos[781] = 90;
				cos[782] = 89;
				cos[783] = 89;
				cos[784] = 88;
				cos[785] = 87;
				cos[786] = 87;
				cos[787] = 86;
				cos[788] = 85;
				cos[789] = 84;
				cos[790] = 84;
				cos[791] = 83;
				cos[792] = 82;
				cos[793] = 82;
				cos[794] = 81;
				cos[795] = 80;
				cos[796] = 80;
				cos[797] = 79;
				cos[798] = 78;
				cos[799] = 78;
				cos[800] = 77;
				cos[801] = 76;
				cos[802] = 76;
				cos[803] = 75;
				cos[804] = 74;
				cos[805] = 74;
				cos[806] = 73;
				cos[807] = 72;
				cos[808] = 72;
				cos[809] = 71;
				cos[810] = 70;
				cos[811] = 70;
				cos[812] = 69;
				cos[813] = 69;
				cos[814] = 68;
				cos[815] = 67;
				cos[816] = 67;
				cos[817] = 66;
				cos[818] = 65;
				cos[819] = 65;
				cos[820] = 64;
				cos[821] = 64;
				cos[822] = 63;
				cos[823] = 62;
				cos[824] = 62;
				cos[825] = 61;
				cos[826] = 61;
				cos[827] = 60;
				cos[828] = 59;
				cos[829] = 59;
				cos[830] = 58;
				cos[831] = 58;
				cos[832] = 57;
				cos[833] = 56;
				cos[834] = 56;
				cos[835] = 55;
				cos[836] = 55;
				cos[837] = 54;
				cos[838] = 54;
				cos[839] = 53;
				cos[840] = 52;
				cos[841] = 52;
				cos[842] = 51;
				cos[843] = 51;
				cos[844] = 50;
				cos[845] = 50;
				cos[846] = 49;
				cos[847] = 49;
				cos[848] = 48;
				cos[849] = 48;
				cos[850] = 47;
				cos[851] = 46;
				cos[852] = 46;
				cos[853] = 45;
				cos[854] = 45;
				cos[855] = 44;
				cos[856] = 44;
				cos[857] = 43;
				cos[858] = 43;
				cos[859] = 42;
				cos[860] = 42;
				cos[861] = 41;
				cos[862] = 41;
				cos[863] = 40;
				cos[864] = 40;
				cos[865] = 39;
				cos[866] = 39;
				cos[867] = 38;
				cos[868] = 38;
				cos[869] = 37;
				cos[870] = 37;
				cos[871] = 36;
				cos[872] = 36;
				cos[873] = 35;
				cos[874] = 35;
				cos[875] = 35;
				cos[876] = 34;
				cos[877] = 34;
				cos[878] = 33;
				cos[879] = 33;
				cos[880] = 32;
				cos[881] = 32;
				cos[882] = 31;
				cos[883] = 31;
				cos[884] = 31;
				cos[885] = 30;
				cos[886] = 30;
				cos[887] = 29;
				cos[888] = 29;
				cos[889] = 28;
				cos[890] = 28;
				cos[891] = 28;
				cos[892] = 27;
				cos[893] = 27;
				cos[894] = 26;
				cos[895] = 26;
				cos[896] = 25;
				cos[897] = 25;
				cos[898] = 25;
				cos[899] = 24;
				cos[900] = 24;
				cos[901] = 24;
				cos[902] = 23;
				cos[903] = 23;
				cos[904] = 22;
				cos[905] = 22;
				cos[906] = 22;
				cos[907] = 21;
				cos[908] = 21;
				cos[909] = 21;
				cos[910] = 20;
				cos[911] = 20;
				cos[912] = 19;
				cos[913] = 19;
				cos[914] = 19;
				cos[915] = 18;
				cos[916] = 18;
				cos[917] = 18;
				cos[918] = 17;
				cos[919] = 17;
				cos[920] = 17;
				cos[921] = 16;
				cos[922] = 16;
				cos[923] = 16;
				cos[924] = 15;
				cos[925] = 15;
				cos[926] = 15;
				cos[927] = 15;
				cos[928] = 14;
				cos[929] = 14;
				cos[930] = 14;
				cos[931] = 13;
				cos[932] = 13;
				cos[933] = 13;
				cos[934] = 12;
				cos[935] = 12;
				cos[936] = 12;
				cos[937] = 12;
				cos[938] = 11;
				cos[939] = 11;
				cos[940] = 11;
				cos[941] = 11;
				cos[942] = 10;
				cos[943] = 10;
				cos[944] = 10;
				cos[945] = 9;
				cos[946] = 9;
				cos[947] = 9;
				cos[948] = 9;
				cos[949] = 8;
				cos[950] = 8;
				cos[951] = 8;
				cos[952] = 8;
				cos[953] = 8;
				cos[954] = 7;
				cos[955] = 7;
				cos[956] = 7;
				cos[957] = 7;
				cos[958] = 6;
				cos[959] = 6;
				cos[960] = 6;
				cos[961] = 6;
				cos[962] = 6;
				cos[963] = 5;
				cos[964] = 5;
				cos[965] = 5;
				cos[966] = 5;
				cos[967] = 5;
				cos[968] = 5;
				cos[969] = 4;
				cos[970] = 4;
				cos[971] = 4;
				cos[972] = 4;
				cos[973] = 4;
				cos[974] = 4;
				cos[975] = 3;
				cos[976] = 3;
				cos[977] = 3;
				cos[978] = 3;
				cos[979] = 3;
				cos[980] = 3;
				cos[981] = 2;
				cos[982] = 2;
				cos[983] = 2;
				cos[984] = 2;
				cos[985] = 2;
				cos[986] = 2;
				cos[987] = 2;
				cos[988] = 2;
				cos[989] = 1;
				cos[990] = 1;
				cos[991] = 1;
				cos[992] = 1;
				cos[993] = 1;
				cos[994] = 1;
				cos[995] = 1;
				cos[996] = 1;
				cos[997] = 1;
				cos[998] = 1;
				cos[999] = 1;
				cos[1000] = 0;
				cos[1001] = 0;
				cos[1002] = 0;
				cos[1003] = 0;
				cos[1004] = 0;
				cos[1005] = 0;
				cos[1006] = 0;
				cos[1007] = 0;
				cos[1008] = 0;
				cos[1009] = 0;
				cos[1010] = 0;
				cos[1011] = 0;
				cos[1012] = 0;
				cos[1013] = 0;
				cos[1014] = 0;
				cos[1015] = 0;
				cos[1016] = 0;
				cos[1017] = 0;
				cos[1018] = 0;
				cos[1019] = 0;
				cos[1020] = 0;
				cos[1021] = 0;
				cos[1022] = 0;
				cos[1023] = 0;
				cos[1024] = 0;
				cos[1025] = 0;
				cos[1026] = 0;
				cos[1027] = 0;
				cos[1028] = 0;
				cos[1029] = 0;
				cos[1030] = 0;
				cos[1031] = 0;
				cos[1032] = 0;
				cos[1033] = 0;
				cos[1034] = 0;
				cos[1035] = 0;
				cos[1036] = 0;
				cos[1037] = 0;
				cos[1038] = 0;
				cos[1039] = 0;
				cos[1040] = 0;
				cos[1041] = 0;
				cos[1042] = 0;
				cos[1043] = 0;
				cos[1044] = 0;
				cos[1045] = 0;
				cos[1046] = 0;
				cos[1047] = 0;
				cos[1048] = 0;
				cos[1049] = 1;
				cos[1050] = 1;
				cos[1051] = 1;
				cos[1052] = 1;
				cos[1053] = 1;
				cos[1054] = 1;
				cos[1055] = 1;
				cos[1056] = 1;
				cos[1057] = 1;
				cos[1058] = 1;
				cos[1059] = 1;
				cos[1060] = 2;
				cos[1061] = 2;
				cos[1062] = 2;
				cos[1063] = 2;
				cos[1064] = 2;
				cos[1065] = 2;
				cos[1066] = 2;
				cos[1067] = 2;
				cos[1068] = 3;
				cos[1069] = 3;
				cos[1070] = 3;
				cos[1071] = 3;
				cos[1072] = 3;
				cos[1073] = 3;
				cos[1074] = 4;
				cos[1075] = 4;
				cos[1076] = 4;
				cos[1077] = 4;
				cos[1078] = 4;
				cos[1079] = 4;
				cos[1080] = 5;
				cos[1081] = 5;
				cos[1082] = 5;
				cos[1083] = 5;
				cos[1084] = 5;
				cos[1085] = 5;
				cos[1086] = 6;
				cos[1087] = 6;
				cos[1088] = 6;
				cos[1089] = 6;
				cos[1090] = 6;
				cos[1091] = 7;
				cos[1092] = 7;
				cos[1093] = 7;
				cos[1094] = 7;
				cos[1095] = 8;
				cos[1096] = 8;
				cos[1097] = 8;
				cos[1098] = 8;
				cos[1099] = 8;
				cos[1100] = 9;
				cos[1101] = 9;
				cos[1102] = 9;
				cos[1103] = 9;
				cos[1104] = 10;
				cos[1105] = 10;
				cos[1106] = 10;
				cos[1107] = 11;
				cos[1108] = 11;
				cos[1109] = 11;
				cos[1110] = 11;
				cos[1111] = 12;
				cos[1112] = 12;
				cos[1113] = 12;
				cos[1114] = 12;
				cos[1115] = 13;
				cos[1116] = 13;
				cos[1117] = 13;
				cos[1118] = 14;
				cos[1119] = 14;
				cos[1120] = 14;
				cos[1121] = 15;
				cos[1122] = 15;
				cos[1123] = 15;
				cos[1124] = 15;
				cos[1125] = 16;
				cos[1126] = 16;
				cos[1127] = 16;
				cos[1128] = 17;
				cos[1129] = 17;
				cos[1130] = 17;
				cos[1131] = 18;
				cos[1132] = 18;
				cos[1133] = 18;
				cos[1134] = 19;
				cos[1135] = 19;
				cos[1136] = 19;
				cos[1137] = 20;
				cos[1138] = 20;
				cos[1139] = 21;
				cos[1140] = 21;
				cos[1141] = 21;
				cos[1142] = 22;
				cos[1143] = 22;
				cos[1144] = 22;
				cos[1145] = 23;
				cos[1146] = 23;
				cos[1147] = 24;
				cos[1148] = 24;
				cos[1149] = 24;
				cos[1150] = 25;
				cos[1151] = 25;
				cos[1152] = 25;
				cos[1153] = 26;
				cos[1154] = 26;
				cos[1155] = 27;
				cos[1156] = 27;
				cos[1157] = 28;
				cos[1158] = 28;
				cos[1159] = 28;
				cos[1160] = 29;
				cos[1161] = 29;
				cos[1162] = 30;
				cos[1163] = 30;
				cos[1164] = 31;
				cos[1165] = 31;
				cos[1166] = 31;
				cos[1167] = 32;
				cos[1168] = 32;
				cos[1169] = 33;
				cos[1170] = 33;
				cos[1171] = 34;
				cos[1172] = 34;
				cos[1173] = 35;
				cos[1174] = 35;
				cos[1175] = 35;
				cos[1176] = 36;
				cos[1177] = 36;
				cos[1178] = 37;
				cos[1179] = 37;
				cos[1180] = 38;
				cos[1181] = 38;
				cos[1182] = 39;
				cos[1183] = 39;
				cos[1184] = 40;
				cos[1185] = 40;
				cos[1186] = 41;
				cos[1187] = 41;
				cos[1188] = 42;
				cos[1189] = 42;
				cos[1190] = 43;
				cos[1191] = 43;
				cos[1192] = 44;
				cos[1193] = 44;
				cos[1194] = 45;
				cos[1195] = 45;
				cos[1196] = 46;
				cos[1197] = 46;
				cos[1198] = 47;
				cos[1199] = 48;
				cos[1200] = 48;
				cos[1201] = 49;
				cos[1202] = 49;
				cos[1203] = 50;
				cos[1204] = 50;
				cos[1205] = 51;
				cos[1206] = 51;
				cos[1207] = 52;
				cos[1208] = 52;
				cos[1209] = 53;
				cos[1210] = 54;
				cos[1211] = 54;
				cos[1212] = 55;
				cos[1213] = 55;
				cos[1214] = 56;
				cos[1215] = 56;
				cos[1216] = 57;
				cos[1217] = 58;
				cos[1218] = 58;
				cos[1219] = 59;
				cos[1220] = 59;
				cos[1221] = 60;
				cos[1222] = 61;
				cos[1223] = 61;
				cos[1224] = 62;
				cos[1225] = 62;
				cos[1226] = 63;
				cos[1227] = 64;
				cos[1228] = 64;
				cos[1229] = 65;
				cos[1230] = 65;
				cos[1231] = 66;
				cos[1232] = 67;
				cos[1233] = 67;
				cos[1234] = 68;
				cos[1235] = 69;
				cos[1236] = 69;
				cos[1237] = 70;
				cos[1238] = 70;
				cos[1239] = 71;
				cos[1240] = 72;
				cos[1241] = 72;
				cos[1242] = 73;
				cos[1243] = 74;
				cos[1244] = 74;
				cos[1245] = 75;
				cos[1246] = 76;
				cos[1247] = 76;
				cos[1248] = 77;
				cos[1249] = 78;
				cos[1250] = 78;
				cos[1251] = 79;
				cos[1252] = 80;
				cos[1253] = 80;
				cos[1254] = 81;
				cos[1255] = 82;
				cos[1256] = 82;
				cos[1257] = 83;
				cos[1258] = 84;
				cos[1259] = 84;
				cos[1260] = 85;
				cos[1261] = 86;
				cos[1262] = 87;
				cos[1263] = 87;
				cos[1264] = 88;
				cos[1265] = 89;
				cos[1266] = 89;
				cos[1267] = 90;
				cos[1268] = 91;
				cos[1269] = 91;
				cos[1270] = 92;
				cos[1271] = 93;
				cos[1272] = 94;
				cos[1273] = 94;
				cos[1274] = 95;
				cos[1275] = 96;
				cos[1276] = 97;
				cos[1277] = 97;
				cos[1278] = 98;
				cos[1279] = 99;
				cos[1280] = 99;
				cos[1281] = 100;
				cos[1282] = 101;
				cos[1283] = 102;
				cos[1284] = 102;
				cos[1285] = 103;
				cos[1286] = 104;
				cos[1287] = 105;
				cos[1288] = 105;
				cos[1289] = 106;
				cos[1290] = 107;
				cos[1291] = 108;
				cos[1292] = 109;
				cos[1293] = 109;
				cos[1294] = 110;
				cos[1295] = 111;
				cos[1296] = 112;
				cos[1297] = 112;
				cos[1298] = 113;
				cos[1299] = 114;
				cos[1300] = 115;
				cos[1301] = 116;
				cos[1302] = 116;
				cos[1303] = 117;
				cos[1304] = 118;
				cos[1305] = 119;
				cos[1306] = 119;
				cos[1307] = 120;
				cos[1308] = 121;
				cos[1309] = 122;
				cos[1310] = 123;
				cos[1311] = 123;
				cos[1312] = 124;
				cos[1313] = 125;
				cos[1314] = 126;
				cos[1315] = 127;
				cos[1316] = 128;
				cos[1317] = 128;
				cos[1318] = 129;
				cos[1319] = 130;
				cos[1320] = 131;
				cos[1321] = 132;
				cos[1322] = 132;
				cos[1323] = 133;
				cos[1324] = 134;
				cos[1325] = 135;
				cos[1326] = 136;
				cos[1327] = 137;
				cos[1328] = 138;
				cos[1329] = 138;
				cos[1330] = 139;
				cos[1331] = 140;
				cos[1332] = 141;
				cos[1333] = 142;
				cos[1334] = 143;
				cos[1335] = 143;
				cos[1336] = 144;
				cos[1337] = 145;
				cos[1338] = 146;
				cos[1339] = 147;
				cos[1340] = 148;
				cos[1341] = 149;
				cos[1342] = 149;
				cos[1343] = 150;
				cos[1344] = 151;
				cos[1345] = 152;
				cos[1346] = 153;
				cos[1347] = 154;
				cos[1348] = 155;
				cos[1349] = 156;
				cos[1350] = 156;
				cos[1351] = 157;
				cos[1352] = 158;
				cos[1353] = 159;
				cos[1354] = 160;
				cos[1355] = 161;
				cos[1356] = 162;
				cos[1357] = 163;
				cos[1358] = 164;
				cos[1359] = 164;
				cos[1360] = 165;
				cos[1361] = 166;
				cos[1362] = 167;
				cos[1363] = 168;
				cos[1364] = 169;
				cos[1365] = 170;
				cos[1366] = 171;
				cos[1367] = 172;
				cos[1368] = 173;
				cos[1369] = 174;
				cos[1370] = 174;
				cos[1371] = 175;
				cos[1372] = 176;
				cos[1373] = 177;
				cos[1374] = 178;
				cos[1375] = 179;
				cos[1376] = 180;
				cos[1377] = 181;
				cos[1378] = 182;
				cos[1379] = 183;
				cos[1380] = 184;
				cos[1381] = 185;
				cos[1382] = 185;
				cos[1383] = 186;
				cos[1384] = 187;
				cos[1385] = 188;
				cos[1386] = 189;
				cos[1387] = 190;
				cos[1388] = 191;
				cos[1389] = 192;
				cos[1390] = 193;
				cos[1391] = 194;
				cos[1392] = 195;
				cos[1393] = 196;
				cos[1394] = 197;
				cos[1395] = 198;
				cos[1396] = 199;
				cos[1397] = 200;
				cos[1398] = 201;
				cos[1399] = 202;
				cos[1400] = 203;
				cos[1401] = 203;
				cos[1402] = 204;
				cos[1403] = 205;
				cos[1404] = 206;
				cos[1405] = 207;
				cos[1406] = 208;
				cos[1407] = 209;
				cos[1408] = 210;
				cos[1409] = 211;
				cos[1410] = 212;
				cos[1411] = 213;
				cos[1412] = 214;
				cos[1413] = 215;
				cos[1414] = 216;
				cos[1415] = 217;
				cos[1416] = 218;
				cos[1417] = 219;
				cos[1418] = 220;
				cos[1419] = 221;
				cos[1420] = 222;
				cos[1421] = 223;
				cos[1422] = 224;
				cos[1423] = 225;
				cos[1424] = 226;
				cos[1425] = 227;
				cos[1426] = 228;
				cos[1427] = 229;
				cos[1428] = 230;
				cos[1429] = 231;
				cos[1430] = 232;
				cos[1431] = 233;
				cos[1432] = 234;
				cos[1433] = 235;
				cos[1434] = 236;
				cos[1435] = 237;
				cos[1436] = 238;
				cos[1437] = 239;
				cos[1438] = 240;
				cos[1439] = 241;
				cos[1440] = 242;
				cos[1441] = 243;
				cos[1442] = 244;
				cos[1443] = 245;
				cos[1444] = 246;
				cos[1445] = 247;
				cos[1446] = 248;
				cos[1447] = 249;
				cos[1448] = 250;
				cos[1449] = 251;
				cos[1450] = 252;
				cos[1451] = 253;
				cos[1452] = 254;
				cos[1453] = 255;
				cos[1454] = 256;
				cos[1455] = 257;
				cos[1456] = 258;
				cos[1457] = 259;
				cos[1458] = 260;
				cos[1459] = 261;
				cos[1460] = 262;
				cos[1461] = 263;
				cos[1462] = 264;
				cos[1463] = 265;
				cos[1464] = 266;
				cos[1465] = 267;
				cos[1466] = 268;
				cos[1467] = 269;
				cos[1468] = 270;
				cos[1469] = 271;
				cos[1470] = 272;
				cos[1471] = 273;
				cos[1472] = 274;
				cos[1473] = 275;
				cos[1474] = 276;
				cos[1475] = 277;
				cos[1476] = 278;
				cos[1477] = 279;
				cos[1478] = 280;
				cos[1479] = 281;
				cos[1480] = 282;
				cos[1481] = 284;
				cos[1482] = 285;
				cos[1483] = 286;
				cos[1484] = 287;
				cos[1485] = 288;
				cos[1486] = 289;
				cos[1487] = 290;
				cos[1488] = 291;
				cos[1489] = 292;
				cos[1490] = 293;
				cos[1491] = 294;
				cos[1492] = 295;
				cos[1493] = 296;
				cos[1494] = 297;
				cos[1495] = 298;
				cos[1496] = 299;
				cos[1497] = 300;
				cos[1498] = 301;
				cos[1499] = 302;
				cos[1500] = 303;
				cos[1501] = 304;
				cos[1502] = 305;
				cos[1503] = 306;
				cos[1504] = 307;
				cos[1505] = 308;
				cos[1506] = 309;
				cos[1507] = 311;
				cos[1508] = 312;
				cos[1509] = 313;
				cos[1510] = 314;
				cos[1511] = 315;
				cos[1512] = 316;
				cos[1513] = 317;
				cos[1514] = 318;
				cos[1515] = 319;
				cos[1516] = 320;
				cos[1517] = 321;
				cos[1518] = 322;
				cos[1519] = 323;
				cos[1520] = 324;
				cos[1521] = 325;
				cos[1522] = 326;
				cos[1523] = 327;
				cos[1524] = 328;
				cos[1525] = 329;
				cos[1526] = 330;
				cos[1527] = 331;
				cos[1528] = 332;
				cos[1529] = 334;
				cos[1530] = 335;
				cos[1531] = 336;
				cos[1532] = 337;
				cos[1533] = 338;
				cos[1534] = 339;
				cos[1535] = 340;
				cos[1536] = 341;
				cos[1537] = 342;
				cos[1538] = 343;
				cos[1539] = 344;
				cos[1540] = 345;
				cos[1541] = 346;
				cos[1542] = 347;
				cos[1543] = 348;
				cos[1544] = 349;
				cos[1545] = 350;
				cos[1546] = 351;
				cos[1547] = 352;
				cos[1548] = 353;
				cos[1549] = 354;
				cos[1550] = 355;
				cos[1551] = 357;
				cos[1552] = 358;
				cos[1553] = 359;
				cos[1554] = 360;
				cos[1555] = 361;
				cos[1556] = 362;
				cos[1557] = 363;
				cos[1558] = 364;
				cos[1559] = 365;
				cos[1560] = 366;
				cos[1561] = 367;
				cos[1562] = 368;
				cos[1563] = 369;
				cos[1564] = 370;
				cos[1565] = 371;
				cos[1566] = 372;
				cos[1567] = 373;
				cos[1568] = 374;
				cos[1569] = 375;
				cos[1570] = 376;
				cos[1571] = 377;
				cos[1572] = 378;
				cos[1573] = 379;
				cos[1574] = 381;
				cos[1575] = 382;
				cos[1576] = 383;
				cos[1577] = 384;
				cos[1578] = 385;
				cos[1579] = 386;
				cos[1580] = 387;
				cos[1581] = 388;
				cos[1582] = 389;
				cos[1583] = 390;
				cos[1584] = 391;
				cos[1585] = 392;
				cos[1586] = 393;
				cos[1587] = 394;
				cos[1588] = 395;
				cos[1589] = 396;
				cos[1590] = 397;
				cos[1591] = 398;
				cos[1592] = 399;
				cos[1593] = 400;
				cos[1594] = 401;
				cos[1595] = 402;
				cos[1596] = 403;
				cos[1597] = 404;
				cos[1598] = 405;
				cos[1599] = 406;
				cos[1600] = 407;
				cos[1601] = 408;
				cos[1602] = 409;
				cos[1603] = 411;
				cos[1604] = 412;
				cos[1605] = 413;
				cos[1606] = 414;
				cos[1607] = 415;
				cos[1608] = 416;
				cos[1609] = 417;
				cos[1610] = 418;
				cos[1611] = 419;
				cos[1612] = 420;
				cos[1613] = 421;
				cos[1614] = 422;
				cos[1615] = 423;
				cos[1616] = 424;
				cos[1617] = 425;
				cos[1618] = 426;
				cos[1619] = 427;
				cos[1620] = 428;
				cos[1621] = 429;
				cos[1622] = 430;
				cos[1623] = 431;
				cos[1624] = 432;
				cos[1625] = 433;
				cos[1626] = 434;
				cos[1627] = 435;
				cos[1628] = 436;
				cos[1629] = 437;
				cos[1630] = 438;
				cos[1631] = 439;
				cos[1632] = 440;
				cos[1633] = 441;
				cos[1634] = 442;
				cos[1635] = 443;
				cos[1636] = 444;
				cos[1637] = 445;
				cos[1638] = 446;
				cos[1639] = 447;
				cos[1640] = 448;
				cos[1641] = 449;
				cos[1642] = 450;
				cos[1643] = 451;
				cos[1644] = 452;
				cos[1645] = 453;
				cos[1646] = 454;
				cos[1647] = 455;
				cos[1648] = 456;
				cos[1649] = 457;
				cos[1650] = 458;
				cos[1651] = 459;
				cos[1652] = 460;
				cos[1653] = 461;
				cos[1654] = 462;
				cos[1655] = 463;
				cos[1656] = 464;
				cos[1657] = 465;
				cos[1658] = 466;
				cos[1659] = 467;
				cos[1660] = 468;
				cos[1661] = 469;
				cos[1662] = 470;
				cos[1663] = 470;
				cos[1664] = 471;
				cos[1665] = 472;
				cos[1666] = 473;
				cos[1667] = 474;
				cos[1668] = 475;
				cos[1669] = 476;
				cos[1670] = 477;
				cos[1671] = 478;
				cos[1672] = 479;
				cos[1673] = 480;
				cos[1674] = 481;
				cos[1675] = 482;
				cos[1676] = 483;
				cos[1677] = 484;
				cos[1678] = 485;
				cos[1679] = 486;
				cos[1680] = 487;
				cos[1681] = 488;
				cos[1682] = 489;
				cos[1683] = 490;
				cos[1684] = 491;
				cos[1685] = 491;
				cos[1686] = 492;
				cos[1687] = 493;
				cos[1688] = 494;
				cos[1689] = 495;
				cos[1690] = 496;
				cos[1691] = 497;
				cos[1692] = 498;
				cos[1693] = 499;
				cos[1694] = 500;
				cos[1695] = 501;
				cos[1696] = 502;
				cos[1697] = 503;
				cos[1698] = 504;
				cos[1699] = 505;
				cos[1700] = 505;
				cos[1701] = 506;
				cos[1702] = 507;
				cos[1703] = 508;
				cos[1704] = 509;
				cos[1705] = 510;
				cos[1706] = 511;
				cos[1707] = 512;
				cos[1708] = 513;
				cos[1709] = 514;
				cos[1710] = 515;
				cos[1711] = 515;
				cos[1712] = 516;
				cos[1713] = 517;
				cos[1714] = 518;
				cos[1715] = 519;
				cos[1716] = 520;
				cos[1717] = 521;
				cos[1718] = 522;
				cos[1719] = 523;
				cos[1720] = 523;
				cos[1721] = 524;
				cos[1722] = 525;
				cos[1723] = 526;
				cos[1724] = 527;
				cos[1725] = 528;
				cos[1726] = 529;
				cos[1727] = 530;
				cos[1728] = 530;
				cos[1729] = 531;
				cos[1730] = 532;
				cos[1731] = 533;
				cos[1732] = 534;
				cos[1733] = 535;
				cos[1734] = 536;
				cos[1735] = 537;
				cos[1736] = 537;
				cos[1737] = 538;
				cos[1738] = 539;
				cos[1739] = 540;
				cos[1740] = 541;
				cos[1741] = 542;
				cos[1742] = 542;
				cos[1743] = 543;
				cos[1744] = 544;
				cos[1745] = 545;
				cos[1746] = 546;
				cos[1747] = 547;
				cos[1748] = 548;
				cos[1749] = 548;
				cos[1750] = 549;
				cos[1751] = 550;
				cos[1752] = 551;
				cos[1753] = 552;
				cos[1754] = 552;
				cos[1755] = 553;
				cos[1756] = 554;
				cos[1757] = 555;
				cos[1758] = 556;
				cos[1759] = 557;
				cos[1760] = 557;
				cos[1761] = 558;
				cos[1762] = 559;
				cos[1763] = 560;
				cos[1764] = 561;
				cos[1765] = 561;
				cos[1766] = 562;
				cos[1767] = 563;
				cos[1768] = 564;
				cos[1769] = 565;
				cos[1770] = 565;
				cos[1771] = 566;
				cos[1772] = 567;
				cos[1773] = 568;
				cos[1774] = 569;
				cos[1775] = 569;
				cos[1776] = 570;
				cos[1777] = 571;
				cos[1778] = 572;
				cos[1779] = 572;
				cos[1780] = 573;
				cos[1781] = 574;
				cos[1782] = 575;
				cos[1783] = 575;
				cos[1784] = 576;
				cos[1785] = 577;
				cos[1786] = 578;
				cos[1787] = 578;
				cos[1788] = 579;
				cos[1789] = 580;
				cos[1790] = 581;
				cos[1791] = 581;
				cos[1792] = 582;
				cos[1793] = 583;
				cos[1794] = 584;
				cos[1795] = 584;
				cos[1796] = 585;
				cos[1797] = 586;
				cos[1798] = 587;
				cos[1799] = 587;
				cos[1800] = 588;
				cos[1801] = 589;
				cos[1802] = 589;
				cos[1803] = 590;
				cos[1804] = 591;
				cos[1805] = 592;
				cos[1806] = 592;
				cos[1807] = 593;
				cos[1808] = 594;
				cos[1809] = 594;
				cos[1810] = 595;
				cos[1811] = 596;
				cos[1812] = 597;
				cos[1813] = 597;
				cos[1814] = 598;
				cos[1815] = 599;
				cos[1816] = 599;
				cos[1817] = 600;
				cos[1818] = 601;
				cos[1819] = 601;
				cos[1820] = 602;
				cos[1821] = 603;
				cos[1822] = 603;
				cos[1823] = 604;
				cos[1824] = 605;
				cos[1825] = 605;
				cos[1826] = 606;
				cos[1827] = 607;
				cos[1828] = 607;
				cos[1829] = 608;
				cos[1830] = 609;
				cos[1831] = 609;
				cos[1832] = 610;
				cos[1833] = 611;
				cos[1834] = 611;
				cos[1835] = 612;
				cos[1836] = 612;
				cos[1837] = 613;
				cos[1838] = 614;
				cos[1839] = 614;
				cos[1840] = 615;
				cos[1841] = 616;
				cos[1842] = 616;
				cos[1843] = 617;
				cos[1844] = 617;
				cos[1845] = 618;
				cos[1846] = 619;
				cos[1847] = 619;
				cos[1848] = 620;
				cos[1849] = 621;
				cos[1850] = 621;
				cos[1851] = 622;
				cos[1852] = 622;
				cos[1853] = 623;
				cos[1854] = 623;
				cos[1855] = 624;
				cos[1856] = 625;
				cos[1857] = 625;
				cos[1858] = 626;
				cos[1859] = 626;
				cos[1860] = 627;
				cos[1861] = 628;
				cos[1862] = 628;
				cos[1863] = 629;
				cos[1864] = 629;
				cos[1865] = 630;
				cos[1866] = 630;
				cos[1867] = 631;
				cos[1868] = 631;
				cos[1869] = 632;
				cos[1870] = 633;
				cos[1871] = 633;
				cos[1872] = 634;
				cos[1873] = 634;
				cos[1874] = 635;
				cos[1875] = 635;
				cos[1876] = 636;
				cos[1877] = 636;
				cos[1878] = 637;
				cos[1879] = 637;
				cos[1880] = 638;
				cos[1881] = 638;
				cos[1882] = 639;
				cos[1883] = 639;
				cos[1884] = 640;
				cos[1885] = 640;
				cos[1886] = 641;
				cos[1887] = 641;
				cos[1888] = 642;
				cos[1889] = 642;
				cos[1890] = 643;
				cos[1891] = 643;
				cos[1892] = 644;
				cos[1893] = 644;
				cos[1894] = 645;
				cos[1895] = 645;
				cos[1896] = 646;
				cos[1897] = 646;
				cos[1898] = 647;
				cos[1899] = 647;
				cos[1900] = 648;
				cos[1901] = 648;
				cos[1902] = 648;
				cos[1903] = 649;
				cos[1904] = 649;
				cos[1905] = 650;
				cos[1906] = 650;
				cos[1907] = 651;
				cos[1908] = 651;
				cos[1909] = 652;
				cos[1910] = 652;
				cos[1911] = 652;
				cos[1912] = 653;
				cos[1913] = 653;
				cos[1914] = 654;
				cos[1915] = 654;
				cos[1916] = 655;
				cos[1917] = 655;
				cos[1918] = 655;
				cos[1919] = 656;
				cos[1920] = 656;
				cos[1921] = 657;
				cos[1922] = 657;
				cos[1923] = 657;
				cos[1924] = 658;
				cos[1925] = 658;
				cos[1926] = 659;
				cos[1927] = 659;
				cos[1928] = 659;
				cos[1929] = 660;
				cos[1930] = 660;
				cos[1931] = 660;
				cos[1932] = 661;
				cos[1933] = 661;
				cos[1934] = 662;
				cos[1935] = 662;
				cos[1936] = 662;
				cos[1937] = 663;
				cos[1938] = 663;
				cos[1939] = 663;
				cos[1940] = 664;
				cos[1941] = 664;
				cos[1942] = 664;
				cos[1943] = 665;
				cos[1944] = 665;
				cos[1945] = 665;
				cos[1946] = 666;
				cos[1947] = 666;
				cos[1948] = 666;
				cos[1949] = 667;
				cos[1950] = 667;
				cos[1951] = 667;
				cos[1952] = 667;
				cos[1953] = 668;
				cos[1954] = 668;
				cos[1955] = 668;
				cos[1956] = 669;
				cos[1957] = 669;
				cos[1958] = 669;
				cos[1959] = 670;
				cos[1960] = 670;
				cos[1961] = 670;
				cos[1962] = 670;
				cos[1963] = 671;
				cos[1964] = 671;
				cos[1965] = 671;
				cos[1966] = 671;
				cos[1967] = 672;
				cos[1968] = 672;
				cos[1969] = 672;
				cos[1970] = 672;
				cos[1971] = 673;
				cos[1972] = 673;
				cos[1973] = 673;
				cos[1974] = 673;
				cos[1975] = 674;
				cos[1976] = 674;
				cos[1977] = 674;
				cos[1978] = 674;
				cos[1979] = 675;
				cos[1980] = 675;
				cos[1981] = 675;
				cos[1982] = 675;
				cos[1983] = 675;
				cos[1984] = 676;
				cos[1985] = 676;
				cos[1986] = 676;
				cos[1987] = 676;
				cos[1988] = 676;
				cos[1989] = 677;
				cos[1990] = 677;
				cos[1991] = 677;
				cos[1992] = 677;
				cos[1993] = 677;
				cos[1994] = 677;
				cos[1995] = 678;
				cos[1996] = 678;
				cos[1997] = 678;
				cos[1998] = 678;
				cos[1999] = 678;
				cos[2000] = 678;
				cos[2001] = 679;
				cos[2002] = 679;
				cos[2003] = 679;
				cos[2004] = 679;
				cos[2005] = 679;
				cos[2006] = 679;
				cos[2007] = 679;
				cos[2008] = 680;
				cos[2009] = 680;
				cos[2010] = 680;
				cos[2011] = 680;
				cos[2012] = 680;
				cos[2013] = 680;
				cos[2014] = 680;
				cos[2015] = 680;
				cos[2016] = 681;
				cos[2017] = 681;
				cos[2018] = 681;
				cos[2019] = 681;
				cos[2020] = 681;
				cos[2021] = 681;
				cos[2022] = 681;
				cos[2023] = 681;
				cos[2024] = 681;
				cos[2025] = 681;
				cos[2026] = 681;
				cos[2027] = 681;
				cos[2028] = 682;
				cos[2029] = 682;
				cos[2030] = 682;
				cos[2031] = 682;
				cos[2032] = 682;
				cos[2033] = 682;
				cos[2034] = 682;
				cos[2035] = 682;
				cos[2036] = 682;
				cos[2037] = 682;
				cos[2038] = 682;
				cos[2039] = 682;
				cos[2040] = 682;
				cos[2041] = 682;
				cos[2042] = 682;
				cos[2043] = 682;
				cos[2044] = 682;
				cos[2045] = 682;
				cos[2046] = 682;
				cos[2047] = 682;   
    end
endmodule
