module sine_output(counter, sine_out);
    input counter;
    output [15:0] sine_out;

    reg [15:0] sine [0:1023];
    initial
        begin
            sine[0] = 0;
            sine[1] = 268;
            sine[2] = 536;
            sine[3] = 804;
            sine[4] = 1072;
            sine[5] = 1340;
            sine[6] = 1608;
            sine[7] = 1875;
            sine[8] = 2143;
            sine[9] = 2411;
            sine[10] = 2679;
            sine[11] = 2946;
            sine[12] = 3214;
            sine[13] = 3481;
            sine[14] = 3748;
            sine[15] = 4015;
            sine[16] = 4282;
            sine[17] = 4549;
            sine[18] = 4815;
            sine[19] = 5081;
            sine[20] = 5348;
            sine[21] = 5614;
            sine[22] = 5879;
            sine[23] = 6145;
            sine[24] = 6410;
            sine[25] = 6675;
            sine[26] = 6940;
            sine[27] = 7205;
            sine[28] = 7469;
            sine[29] = 7733;
            sine[30] = 7997;
            sine[31] = 8260;
            sine[32] = 8523;
            sine[33] = 8786;
            sine[34] = 9048;
            sine[35] = 9310;
            sine[36] = 9572;
            sine[37] = 9833;
            sine[38] = 10094;
            sine[39] = 10355;
            sine[40] = 10615;
            sine[41] = 10875;
            sine[42] = 11135;
            sine[43] = 11394;
            sine[44] = 11652;
            sine[45] = 11910;
            sine[46] = 12168;
            sine[47] = 12425;
            sine[48] = 12682;
            sine[49] = 12938;
            sine[50] = 13194;
            sine[51] = 13449;
            sine[52] = 13704;
            sine[53] = 13959;
            sine[54] = 14212;
            sine[55] = 14466;
            sine[56] = 14718;
            sine[57] = 14970;
            sine[58] = 15222;
            sine[59] = 15473;
            sine[60] = 15723;
            sine[61] = 15973;
            sine[62] = 16222;
            sine[63] = 16471;
            sine[64] = 16719;
            sine[65] = 16966;
            sine[66] = 17213;
            sine[67] = 17459;
            sine[68] = 17704;
            sine[69] = 17949;
            sine[70] = 18193;
            sine[71] = 18437;
            sine[72] = 18679;
            sine[73] = 18921;
            sine[74] = 19163;
            sine[75] = 19403;
            sine[76] = 19643;
            sine[77] = 19882;
            sine[78] = 20120;
            sine[79] = 20358;
            sine[80] = 20595;
            sine[81] = 20831;
            sine[82] = 21066;
            sine[83] = 21301;
            sine[84] = 21534;
            sine[85] = 21767;
            sine[86] = 21999;
            sine[87] = 22230;
            sine[88] = 22461;
            sine[89] = 22690;
            sine[90] = 22919;
            sine[91] = 23147;
            sine[92] = 23374;
            sine[93] = 23600;
            sine[94] = 23825;
            sine[95] = 24049;
            sine[96] = 24272;
            sine[97] = 24495;
            sine[98] = 24716;
            sine[99] = 24937;
            sine[100] = 25157;
            sine[101] = 25375;
            sine[102] = 25593;
            sine[103] = 25810;
            sine[104] = 26026;
            sine[105] = 26240;
            sine[106] = 26454;
            sine[107] = 26667;
            sine[108] = 26879;
            sine[109] = 27090;
            sine[110] = 27300;
            sine[111] = 27508;
            sine[112] = 27716;
            sine[113] = 27923;
            sine[114] = 28129;
            sine[115] = 28333;
            sine[116] = 28537;
            sine[117] = 28739;
            sine[118] = 28940;
            sine[119] = 29141;
            sine[120] = 29340;
            sine[121] = 29538;
            sine[122] = 29735;
            sine[123] = 29931;
            sine[124] = 30126;
            sine[125] = 30319;
            sine[126] = 30512;
            sine[127] = 30703;
            sine[128] = 30893;
            sine[129] = 31082;
            sine[130] = 31270;
            sine[131] = 31456;
            sine[132] = 31642;
            sine[133] = 31826;
            sine[134] = 32009;
            sine[135] = 32191;
            sine[136] = 32372;
            sine[137] = 32551;
            sine[138] = 32729;
            sine[139] = 32906;
            sine[140] = 33082;
            sine[141] = 33256;
            sine[142] = 33430;
            sine[143] = 33602;
            sine[144] = 33772;
            sine[145] = 33942;
            sine[146] = 34110;
            sine[147] = 34277;
            sine[148] = 34442;
            sine[149] = 34607;
            sine[150] = 34770;
            sine[151] = 34931;
            sine[152] = 35092;
            sine[153] = 35251;
            sine[154] = 35408;
            sine[155] = 35565;
            sine[156] = 35720;
            sine[157] = 35873;
            sine[158] = 36026;
            sine[159] = 36177;
            sine[160] = 36326;
            sine[161] = 36475;
            sine[162] = 36622;
            sine[163] = 36767;
            sine[164] = 36911;
            sine[165] = 37054;
            sine[166] = 37195;
            sine[167] = 37335;
            sine[168] = 37474;
            sine[169] = 37611;
            sine[170] = 37746;
            sine[171] = 37881;
            sine[172] = 38014;
            sine[173] = 38145;
            sine[174] = 38275;
            sine[175] = 38404;
            sine[176] = 38531;
            sine[177] = 38656;
            sine[178] = 38780;
            sine[179] = 38903;
            sine[180] = 39024;
            sine[181] = 39144;
            sine[182] = 39263;
            sine[183] = 39379;
            sine[184] = 39495;
            sine[185] = 39609;
            sine[186] = 39721;
            sine[187] = 39832;
            sine[188] = 39941;
            sine[189] = 40049;
            sine[190] = 40156;
            sine[191] = 40260;
            sine[192] = 40364;
            sine[193] = 40466;
            sine[194] = 40566;
            sine[195] = 40665;
            sine[196] = 40762;
            sine[197] = 40858;
            sine[198] = 40952;
            sine[199] = 41044;
            sine[200] = 41136;
            sine[201] = 41225;
            sine[202] = 41313;
            sine[203] = 41400;
            sine[204] = 41484;
            sine[205] = 41568;
            sine[206] = 41649;
            sine[207] = 41730;
            sine[208] = 41808;
            sine[209] = 41885;
            sine[210] = 41961;
            sine[211] = 42035;
            sine[212] = 42107;
            sine[213] = 42178;
            sine[214] = 42247;
            sine[215] = 42314;
            sine[216] = 42380;
            sine[217] = 42445;
            sine[218] = 42507;
            sine[219] = 42568;
            sine[220] = 42628;
            sine[221] = 42686;
            sine[222] = 42742;
            sine[223] = 42797;
            sine[224] = 42850;
            sine[225] = 42902;
            sine[226] = 42951;
            sine[227] = 43000;
            sine[228] = 43046;
            sine[229] = 43091;
            sine[230] = 43135;
            sine[231] = 43176;
            sine[232] = 43217;
            sine[233] = 43255;
            sine[234] = 43292;
            sine[235] = 43327;
            sine[236] = 43361;
            sine[237] = 43393;
            sine[238] = 43423;
            sine[239] = 43452;
            sine[240] = 43479;
            sine[241] = 43505;
            sine[242] = 43528;
            sine[243] = 43551;
            sine[244] = 43571;
            sine[245] = 43590;
            sine[246] = 43607;
            sine[247] = 43623;
            sine[248] = 43637;
            sine[249] = 43649;
            sine[250] = 43660;
            sine[251] = 43669;
            sine[252] = 43676;
            sine[253] = 43682;
            sine[254] = 43686;
            sine[255] = 43689;
            sine[256] = 43690;
            sine[257] = 43689;
            sine[258] = 43686;
            sine[259] = 43682;
            sine[260] = 43676;
            sine[261] = 43669;
            sine[262] = 43660;
            sine[263] = 43649;
            sine[264] = 43637;
            sine[265] = 43623;
            sine[266] = 43607;
            sine[267] = 43590;
            sine[268] = 43571;
            sine[269] = 43551;
            sine[270] = 43528;
            sine[271] = 43505;
            sine[272] = 43479;
            sine[273] = 43452;
            sine[274] = 43423;
            sine[275] = 43393;
            sine[276] = 43361;
            sine[277] = 43327;
            sine[278] = 43292;
            sine[279] = 43255;
            sine[280] = 43217;
            sine[281] = 43176;
            sine[282] = 43135;
            sine[283] = 43091;
            sine[284] = 43046;
            sine[285] = 43000;
            sine[286] = 42951;
            sine[287] = 42902;
            sine[288] = 42850;
            sine[289] = 42797;
            sine[290] = 42742;
            sine[291] = 42686;
            sine[292] = 42628;
            sine[293] = 42568;
            sine[294] = 42507;
            sine[295] = 42445;
            sine[296] = 42380;
            sine[297] = 42314;
            sine[298] = 42247;
            sine[299] = 42178;
            sine[300] = 42107;
            sine[301] = 42035;
            sine[302] = 41961;
            sine[303] = 41885;
            sine[304] = 41808;
            sine[305] = 41730;
            sine[306] = 41649;
            sine[307] = 41568;
            sine[308] = 41484;
            sine[309] = 41400;
            sine[310] = 41313;
            sine[311] = 41225;
            sine[312] = 41136;
            sine[313] = 41044;
            sine[314] = 40952;
            sine[315] = 40858;
            sine[316] = 40762;
            sine[317] = 40665;
            sine[318] = 40566;
            sine[319] = 40466;
            sine[320] = 40364;
            sine[321] = 40260;
            sine[322] = 40156;
            sine[323] = 40049;
            sine[324] = 39941;
            sine[325] = 39832;
            sine[326] = 39721;
            sine[327] = 39609;
            sine[328] = 39495;
            sine[329] = 39379;
            sine[330] = 39263;
            sine[331] = 39144;
            sine[332] = 39024;
            sine[333] = 38903;
            sine[334] = 38780;
            sine[335] = 38656;
            sine[336] = 38531;
            sine[337] = 38404;
            sine[338] = 38275;
            sine[339] = 38145;
            sine[340] = 38014;
            sine[341] = 37881;
            sine[342] = 37746;
            sine[343] = 37611;
            sine[344] = 37474;
            sine[345] = 37335;
            sine[346] = 37195;
            sine[347] = 37054;
            sine[348] = 36911;
            sine[349] = 36767;
            sine[350] = 36622;
            sine[351] = 36475;
            sine[352] = 36326;
            sine[353] = 36177;
            sine[354] = 36026;
            sine[355] = 35873;
            sine[356] = 35720;
            sine[357] = 35565;
            sine[358] = 35408;
            sine[359] = 35251;
            sine[360] = 35092;
            sine[361] = 34931;
            sine[362] = 34770;
            sine[363] = 34607;
            sine[364] = 34442;
            sine[365] = 34277;
            sine[366] = 34110;
            sine[367] = 33942;
            sine[368] = 33772;
            sine[369] = 33602;
            sine[370] = 33430;
            sine[371] = 33256;
            sine[372] = 33082;
            sine[373] = 32906;
            sine[374] = 32729;
            sine[375] = 32551;
            sine[376] = 32372;
            sine[377] = 32191;
            sine[378] = 32009;
            sine[379] = 31826;
            sine[380] = 31642;
            sine[381] = 31456;
            sine[382] = 31270;
            sine[383] = 31082;
            sine[384] = 30893;
            sine[385] = 30703;
            sine[386] = 30512;
            sine[387] = 30319;
            sine[388] = 30126;
            sine[389] = 29931;
            sine[390] = 29735;
            sine[391] = 29538;
            sine[392] = 29340;
            sine[393] = 29141;
            sine[394] = 28940;
            sine[395] = 28739;
            sine[396] = 28537;
            sine[397] = 28333;
            sine[398] = 28129;
            sine[399] = 27923;
            sine[400] = 27716;
            sine[401] = 27508;
            sine[402] = 27300;
            sine[403] = 27090;
            sine[404] = 26879;
            sine[405] = 26667;
            sine[406] = 26454;
            sine[407] = 26240;
            sine[408] = 26026;
            sine[409] = 25810;
            sine[410] = 25593;
            sine[411] = 25375;
            sine[412] = 25157;
            sine[413] = 24937;
            sine[414] = 24716;
            sine[415] = 24495;
            sine[416] = 24272;
            sine[417] = 24049;
            sine[418] = 23825;
            sine[419] = 23600;
            sine[420] = 23374;
            sine[421] = 23147;
            sine[422] = 22919;
            sine[423] = 22690;
            sine[424] = 22461;
            sine[425] = 22230;
            sine[426] = 21999;
            sine[427] = 21767;
            sine[428] = 21534;
            sine[429] = 21301;
            sine[430] = 21066;
            sine[431] = 20831;
            sine[432] = 20595;
            sine[433] = 20358;
            sine[434] = 20120;
            sine[435] = 19882;
            sine[436] = 19643;
            sine[437] = 19403;
            sine[438] = 19163;
            sine[439] = 18921;
            sine[440] = 18679;
            sine[441] = 18437;
            sine[442] = 18193;
            sine[443] = 17949;
            sine[444] = 17704;
            sine[445] = 17459;
            sine[446] = 17213;
            sine[447] = 16966;
            sine[448] = 16719;
            sine[449] = 16471;
            sine[450] = 16222;
            sine[451] = 15973;
            sine[452] = 15723;
            sine[453] = 15473;
            sine[454] = 15222;
            sine[455] = 14970;
            sine[456] = 14718;
            sine[457] = 14466;
            sine[458] = 14212;
            sine[459] = 13959;
            sine[460] = 13704;
            sine[461] = 13449;
            sine[462] = 13194;
            sine[463] = 12938;
            sine[464] = 12682;
            sine[465] = 12425;
            sine[466] = 12168;
            sine[467] = 11910;
            sine[468] = 11652;
            sine[469] = 11394;
            sine[470] = 11135;
            sine[471] = 10875;
            sine[472] = 10615;
            sine[473] = 10355;
            sine[474] = 10094;
            sine[475] = 9833;
            sine[476] = 9572;
            sine[477] = 9310;
            sine[478] = 9048;
            sine[479] = 8786;
            sine[480] = 8523;
            sine[481] = 8260;
            sine[482] = 7997;
            sine[483] = 7733;
            sine[484] = 7469;
            sine[485] = 7205;
            sine[486] = 6940;
            sine[487] = 6675;
            sine[488] = 6410;
            sine[489] = 6145;
            sine[490] = 5879;
            sine[491] = 5614;
            sine[492] = 5348;
            sine[493] = 5081;
            sine[494] = 4815;
            sine[495] = 4549;
            sine[496] = 4282;
            sine[497] = 4015;
            sine[498] = 3748;
            sine[499] = 3481;
            sine[500] = 3214;
            sine[501] = 2946;
            sine[502] = 2679;
            sine[503] = 2411;
            sine[504] = 2143;
            sine[505] = 1875;
            sine[506] = 1608;
            sine[507] = 1340;
            sine[508] = 1072;
            sine[509] = 804;
            sine[510] = 536;
            sine[511] = 268;
            sine[512] = 0;
            sine[513] = -268;
            sine[514] = -536;
            sine[515] = -804;
            sine[516] = -1072;
            sine[517] = -1340;
            sine[518] = -1608;
            sine[519] = -1875;
            sine[520] = -2143;
            sine[521] = -2411;
            sine[522] = -2679;
            sine[523] = -2946;
            sine[524] = -3214;
            sine[525] = -3481;
            sine[526] = -3748;
            sine[527] = -4015;
            sine[528] = -4282;
            sine[529] = -4549;
            sine[530] = -4815;
            sine[531] = -5081;
            sine[532] = -5348;
            sine[533] = -5614;
            sine[534] = -5879;
            sine[535] = -6145;
            sine[536] = -6410;
            sine[537] = -6675;
            sine[538] = -6940;
            sine[539] = -7205;
            sine[540] = -7469;
            sine[541] = -7733;
            sine[542] = -7997;
            sine[543] = -8260;
            sine[544] = -8523;
            sine[545] = -8786;
            sine[546] = -9048;
            sine[547] = -9310;
            sine[548] = -9572;
            sine[549] = -9833;
            sine[550] = -10094;
            sine[551] = -10355;
            sine[552] = -10615;
            sine[553] = -10875;
            sine[554] = -11135;
            sine[555] = -11394;
            sine[556] = -11652;
            sine[557] = -11910;
            sine[558] = -12168;
            sine[559] = -12425;
            sine[560] = -12682;
            sine[561] = -12938;
            sine[562] = -13194;
            sine[563] = -13449;
            sine[564] = -13704;
            sine[565] = -13959;
            sine[566] = -14212;
            sine[567] = -14466;
            sine[568] = -14718;
            sine[569] = -14970;
            sine[570] = -15222;
            sine[571] = -15473;
            sine[572] = -15723;
            sine[573] = -15973;
            sine[574] = -16222;
            sine[575] = -16471;
            sine[576] = -16719;
            sine[577] = -16966;
            sine[578] = -17213;
            sine[579] = -17459;
            sine[580] = -17704;
            sine[581] = -17949;
            sine[582] = -18193;
            sine[583] = -18437;
            sine[584] = -18679;
            sine[585] = -18921;
            sine[586] = -19163;
            sine[587] = -19403;
            sine[588] = -19643;
            sine[589] = -19882;
            sine[590] = -20120;
            sine[591] = -20358;
            sine[592] = -20595;
            sine[593] = -20831;
            sine[594] = -21066;
            sine[595] = -21301;
            sine[596] = -21534;
            sine[597] = -21767;
            sine[598] = -21999;
            sine[599] = -22230;
            sine[600] = -22461;
            sine[601] = -22690;
            sine[602] = -22919;
            sine[603] = -23147;
            sine[604] = -23374;
            sine[605] = -23600;
            sine[606] = -23825;
            sine[607] = -24049;
            sine[608] = -24272;
            sine[609] = -24495;
            sine[610] = -24716;
            sine[611] = -24937;
            sine[612] = -25157;
            sine[613] = -25375;
            sine[614] = -25593;
            sine[615] = -25810;
            sine[616] = -26026;
            sine[617] = -26240;
            sine[618] = -26454;
            sine[619] = -26667;
            sine[620] = -26879;
            sine[621] = -27090;
            sine[622] = -27300;
            sine[623] = -27508;
            sine[624] = -27716;
            sine[625] = -27923;
            sine[626] = -28129;
            sine[627] = -28333;
            sine[628] = -28537;
            sine[629] = -28739;
            sine[630] = -28940;
            sine[631] = -29141;
            sine[632] = -29340;
            sine[633] = -29538;
            sine[634] = -29735;
            sine[635] = -29931;
            sine[636] = -30126;
            sine[637] = -30319;
            sine[638] = -30512;
            sine[639] = -30703;
            sine[640] = -30893;
            sine[641] = -31082;
            sine[642] = -31270;
            sine[643] = -31456;
            sine[644] = -31642;
            sine[645] = -31826;
            sine[646] = -32009;
            sine[647] = -32191;
            sine[648] = -32372;
            sine[649] = -32551;
            sine[650] = -32729;
            sine[651] = -32906;
            sine[652] = -33082;
            sine[653] = -33256;
            sine[654] = -33430;
            sine[655] = -33602;
            sine[656] = -33772;
            sine[657] = -33942;
            sine[658] = -34110;
            sine[659] = -34277;
            sine[660] = -34442;
            sine[661] = -34607;
            sine[662] = -34770;
            sine[663] = -34931;
            sine[664] = -35092;
            sine[665] = -35251;
            sine[666] = -35408;
            sine[667] = -35565;
            sine[668] = -35720;
            sine[669] = -35873;
            sine[670] = -36026;
            sine[671] = -36177;
            sine[672] = -36326;
            sine[673] = -36475;
            sine[674] = -36622;
            sine[675] = -36767;
            sine[676] = -36911;
            sine[677] = -37054;
            sine[678] = -37195;
            sine[679] = -37335;
            sine[680] = -37474;
            sine[681] = -37611;
            sine[682] = -37746;
            sine[683] = -37881;
            sine[684] = -38014;
            sine[685] = -38145;
            sine[686] = -38275;
            sine[687] = -38404;
            sine[688] = -38531;
            sine[689] = -38656;
            sine[690] = -38780;
            sine[691] = -38903;
            sine[692] = -39024;
            sine[693] = -39144;
            sine[694] = -39263;
            sine[695] = -39379;
            sine[696] = -39495;
            sine[697] = -39609;
            sine[698] = -39721;
            sine[699] = -39832;
            sine[700] = -39941;
            sine[701] = -40049;
            sine[702] = -40156;
            sine[703] = -40260;
            sine[704] = -40364;
            sine[705] = -40466;
            sine[706] = -40566;
            sine[707] = -40665;
            sine[708] = -40762;
            sine[709] = -40858;
            sine[710] = -40952;
            sine[711] = -41044;
            sine[712] = -41136;
            sine[713] = -41225;
            sine[714] = -41313;
            sine[715] = -41400;
            sine[716] = -41484;
            sine[717] = -41568;
            sine[718] = -41649;
            sine[719] = -41730;
            sine[720] = -41808;
            sine[721] = -41885;
            sine[722] = -41961;
            sine[723] = -42035;
            sine[724] = -42107;
            sine[725] = -42178;
            sine[726] = -42247;
            sine[727] = -42314;
            sine[728] = -42380;
            sine[729] = -42445;
            sine[730] = -42507;
            sine[731] = -42568;
            sine[732] = -42628;
            sine[733] = -42686;
            sine[734] = -42742;
            sine[735] = -42797;
            sine[736] = -42850;
            sine[737] = -42902;
            sine[738] = -42951;
            sine[739] = -43000;
            sine[740] = -43046;
            sine[741] = -43091;
            sine[742] = -43135;
            sine[743] = -43176;
            sine[744] = -43217;
            sine[745] = -43255;
            sine[746] = -43292;
            sine[747] = -43327;
            sine[748] = -43361;
            sine[749] = -43393;
            sine[750] = -43423;
            sine[751] = -43452;
            sine[752] = -43479;
            sine[753] = -43505;
            sine[754] = -43528;
            sine[755] = -43551;
            sine[756] = -43571;
            sine[757] = -43590;
            sine[758] = -43607;
            sine[759] = -43623;
            sine[760] = -43637;
            sine[761] = -43649;
            sine[762] = -43660;
            sine[763] = -43669;
            sine[764] = -43676;
            sine[765] = -43682;
            sine[766] = -43686;
            sine[767] = -43689;
            sine[768] = -43690;
            sine[769] = -43689;
            sine[770] = -43686;
            sine[771] = -43682;
            sine[772] = -43676;
            sine[773] = -43669;
            sine[774] = -43660;
            sine[775] = -43649;
            sine[776] = -43637;
            sine[777] = -43623;
            sine[778] = -43607;
            sine[779] = -43590;
            sine[780] = -43571;
            sine[781] = -43551;
            sine[782] = -43528;
            sine[783] = -43505;
            sine[784] = -43479;
            sine[785] = -43452;
            sine[786] = -43423;
            sine[787] = -43393;
            sine[788] = -43361;
            sine[789] = -43327;
            sine[790] = -43292;
            sine[791] = -43255;
            sine[792] = -43217;
            sine[793] = -43176;
            sine[794] = -43135;
            sine[795] = -43091;
            sine[796] = -43046;
            sine[797] = -43000;
            sine[798] = -42951;
            sine[799] = -42902;
            sine[800] = -42850;
            sine[801] = -42797;
            sine[802] = -42742;
            sine[803] = -42686;
            sine[804] = -42628;
            sine[805] = -42568;
            sine[806] = -42507;
            sine[807] = -42445;
            sine[808] = -42380;
            sine[809] = -42314;
            sine[810] = -42247;
            sine[811] = -42178;
            sine[812] = -42107;
            sine[813] = -42035;
            sine[814] = -41961;
            sine[815] = -41885;
            sine[816] = -41808;
            sine[817] = -41730;
            sine[818] = -41649;
            sine[819] = -41568;
            sine[820] = -41484;
            sine[821] = -41400;
            sine[822] = -41313;
            sine[823] = -41225;
            sine[824] = -41136;
            sine[825] = -41044;
            sine[826] = -40952;
            sine[827] = -40858;
            sine[828] = -40762;
            sine[829] = -40665;
            sine[830] = -40566;
            sine[831] = -40466;
            sine[832] = -40364;
            sine[833] = -40260;
            sine[834] = -40156;
            sine[835] = -40049;
            sine[836] = -39941;
            sine[837] = -39832;
            sine[838] = -39721;
            sine[839] = -39609;
            sine[840] = -39495;
            sine[841] = -39379;
            sine[842] = -39263;
            sine[843] = -39144;
            sine[844] = -39024;
            sine[845] = -38903;
            sine[846] = -38780;
            sine[847] = -38656;
            sine[848] = -38531;
            sine[849] = -38404;
            sine[850] = -38275;
            sine[851] = -38145;
            sine[852] = -38014;
            sine[853] = -37881;
            sine[854] = -37746;
            sine[855] = -37611;
            sine[856] = -37474;
            sine[857] = -37335;
            sine[858] = -37195;
            sine[859] = -37054;
            sine[860] = -36911;
            sine[861] = -36767;
            sine[862] = -36622;
            sine[863] = -36475;
            sine[864] = -36326;
            sine[865] = -36177;
            sine[866] = -36026;
            sine[867] = -35873;
            sine[868] = -35720;
            sine[869] = -35565;
            sine[870] = -35408;
            sine[871] = -35251;
            sine[872] = -35092;
            sine[873] = -34931;
            sine[874] = -34770;
            sine[875] = -34607;
            sine[876] = -34442;
            sine[877] = -34277;
            sine[878] = -34110;
            sine[879] = -33942;
            sine[880] = -33772;
            sine[881] = -33602;
            sine[882] = -33430;
            sine[883] = -33256;
            sine[884] = -33082;
            sine[885] = -32906;
            sine[886] = -32729;
            sine[887] = -32551;
            sine[888] = -32372;
            sine[889] = -32191;
            sine[890] = -32009;
            sine[891] = -31826;
            sine[892] = -31642;
            sine[893] = -31456;
            sine[894] = -31270;
            sine[895] = -31082;
            sine[896] = -30893;
            sine[897] = -30703;
            sine[898] = -30512;
            sine[899] = -30319;
            sine[900] = -30126;
            sine[901] = -29931;
            sine[902] = -29735;
            sine[903] = -29538;
            sine[904] = -29340;
            sine[905] = -29141;
            sine[906] = -28940;
            sine[907] = -28739;
            sine[908] = -28537;
            sine[909] = -28333;
            sine[910] = -28129;
            sine[911] = -27923;
            sine[912] = -27716;
            sine[913] = -27508;
            sine[914] = -27300;
            sine[915] = -27090;
            sine[916] = -26879;
            sine[917] = -26667;
            sine[918] = -26454;
            sine[919] = -26240;
            sine[920] = -26026;
            sine[921] = -25810;
            sine[922] = -25593;
            sine[923] = -25375;
            sine[924] = -25157;
            sine[925] = -24937;
            sine[926] = -24716;
            sine[927] = -24495;
            sine[928] = -24272;
            sine[929] = -24049;
            sine[930] = -23825;
            sine[931] = -23600;
            sine[932] = -23374;
            sine[933] = -23147;
            sine[934] = -22919;
            sine[935] = -22690;
            sine[936] = -22461;
            sine[937] = -22230;
            sine[938] = -21999;
            sine[939] = -21767;
            sine[940] = -21534;
            sine[941] = -21301;
            sine[942] = -21066;
            sine[943] = -20831;
            sine[944] = -20595;
            sine[945] = -20358;
            sine[946] = -20120;
            sine[947] = -19882;
            sine[948] = -19643;
            sine[949] = -19403;
            sine[950] = -19163;
            sine[951] = -18921;
            sine[952] = -18679;
            sine[953] = -18437;
            sine[954] = -18193;
            sine[955] = -17949;
            sine[956] = -17704;
            sine[957] = -17459;
            sine[958] = -17213;
            sine[959] = -16966;
            sine[960] = -16719;
            sine[961] = -16471;
            sine[962] = -16222;
            sine[963] = -15973;
            sine[964] = -15723;
            sine[965] = -15473;
            sine[966] = -15222;
            sine[967] = -14970;
            sine[968] = -14718;
            sine[969] = -14466;
            sine[970] = -14212;
            sine[971] = -13959;
            sine[972] = -13704;
            sine[973] = -13449;
            sine[974] = -13194;
            sine[975] = -12938;
            sine[976] = -12682;
            sine[977] = -12425;
            sine[978] = -12168;
            sine[979] = -11910;
            sine[980] = -11652;
            sine[981] = -11394;
            sine[982] = -11135;
            sine[983] = -10875;
            sine[984] = -10615;
            sine[985] = -10355;
            sine[986] = -10094;
            sine[987] = -9833;
            sine[988] = -9572;
            sine[989] = -9310;
            sine[990] = -9048;
            sine[991] = -8786;
            sine[992] = -8523;
            sine[993] = -8260;
            sine[994] = -7997;
            sine[995] = -7733;
            sine[996] = -7469;
            sine[997] = -7205;
            sine[998] = -6940;
            sine[999] = -6675;
            sine[1000] = -6410;
            sine[1001] = -6145;
            sine[1002] = -5879;
            sine[1003] = -5614;
            sine[1004] = -5348;
            sine[1005] = -5081;
            sine[1006] = -4815;
            sine[1007] = -4549;
            sine[1008] = -4282;
            sine[1009] = -4015;
            sine[1010] = -3748;
            sine[1011] = -3481;
            sine[1012] = -3214;
            sine[1013] = -2946;
            sine[1014] = -2679;
            sine[1015] = -2411;
            sine[1016] = -2143;
            sine[1017] = -1875;
            sine[1018] = -1608;
            sine[1019] = -1340;
            sine[1020] = -1072;
            sine[1021] = -804;
            sine[1022] = -536;
            sine[1023] = -268;
        end
    assign sine_out = sine[counter];
endmodule
