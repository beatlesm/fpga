module changevalue (
	output fp_gpio<0>
);

assign fp_gpio<0> = 1'b1;
endmodule
