module changevalue (PPS_IN_INT);

output PPS_IN_INT;
PPS_IN_INT <= 1;

endmodule


