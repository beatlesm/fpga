module input_signal_adv(radio_clk, codeword1, codeword2, get_tx);
   input radio_clk;
   input [31:0] codeword1;
   input [31:0] codeword2;


   output [31:0] get_tx;
   reg [31:0] phase_acc1;
   reg [31:0] phase_acc2;
   reg [31:0] tx_out;

/*   
   always @(posedge radio_clk) begin
        if (count == 0) begin
            codeword = 920030940;
        end
        if (codeword_ch) begin
            count = count + 1;
            codeword = codeword_sr;
        end
    end*/
   // Square Wave
  /* 
   always @(posedge radio_clk) begin
      counter = counter + 1;
      if (counter[1] == 1) begin
      	tx_out[31:16] <= 16'b1010101010101010;
      	tx_out[15:0] <= 16'b1010101010101010;
	end 
      else begin
      	tx_out[31:16] <= 16'b0000000000000000;
      	tx_out[15:0] <= 16'b0000000000000000;
	end
   end
*/
    always @(posedge radio_clk) begin
        phase_acc1 = phase_acc1 + codeword1;
		phase_acc2 = phase_acc2 + codeword2;
        tx_out[10:0] = sine[phase_acc1[31:21]] + sine[phase_acc2[31:21]];
        tx_out[31:11] = 21'b000000000000000000000;
    end
   assign get_tx = tx_out;


// SINE LOOKUP TABLE
    reg [9:0] sine [0:2047];
    initial
        begin
                sine[0] = 341;
                sine[1] = 342;
                sine[2] = 343;
                sine[3] = 344;
                sine[4] = 345;
                sine[5] = 346;
                sine[6] = 347;
                sine[7] = 348;
                sine[8] = 349;
                sine[9] = 350;
                sine[10] = 351;
                sine[11] = 352;
                sine[12] = 353;
                sine[13] = 354;
                sine[14] = 355;
                sine[15] = 356;
                sine[16] = 357;
                sine[17] = 358;
                sine[18] = 359;
                sine[19] = 360;
                sine[20] = 361;
                sine[21] = 362;
                sine[22] = 363;
                sine[23] = 365;
                sine[24] = 366;
                sine[25] = 367;
                sine[26] = 368;
                sine[27] = 369;
                sine[28] = 370;
                sine[29] = 371;
                sine[30] = 372;
                sine[31] = 373;
                sine[32] = 374;
                sine[33] = 375;
                sine[34] = 376;
                sine[35] = 377;
                sine[36] = 378;
                sine[37] = 379;
                sine[38] = 380;
                sine[39] = 381;
                sine[40] = 382;
                sine[41] = 383;
                sine[42] = 384;
                sine[43] = 385;
                sine[44] = 386;
                sine[45] = 387;
                sine[46] = 388;
                sine[47] = 390;
                sine[48] = 391;
                sine[49] = 392;
                sine[50] = 393;
                sine[51] = 394;
                sine[52] = 395;
                sine[53] = 396;
                sine[54] = 397;
                sine[55] = 398;
                sine[56] = 399;
                sine[57] = 400;
                sine[58] = 401;
                sine[59] = 402;
                sine[60] = 403;
                sine[61] = 404;
                sine[62] = 405;
                sine[63] = 406;
                sine[64] = 407;
                sine[65] = 408;
                sine[66] = 409;
                sine[67] = 410;
                sine[68] = 411;
                sine[69] = 412;
                sine[70] = 413;
                sine[71] = 414;
                sine[72] = 415;
                sine[73] = 416;
                sine[74] = 417;
                sine[75] = 418;
                sine[76] = 419;
                sine[77] = 420;
                sine[78] = 421;
                sine[79] = 422;
                sine[80] = 423;
                sine[81] = 424;
                sine[82] = 425;
                sine[83] = 426;
                sine[84] = 427;
                sine[85] = 428;
                sine[86] = 429;
                sine[87] = 430;
                sine[88] = 431;
                sine[89] = 432;
                sine[90] = 433;
                sine[91] = 434;
                sine[92] = 435;
                sine[93] = 436;
                sine[94] = 437;
                sine[95] = 438;
                sine[96] = 439;
                sine[97] = 440;
                sine[98] = 441;
                sine[99] = 442;
                sine[100] = 443;
                sine[101] = 444;
                sine[102] = 445;
                sine[103] = 446;
                sine[104] = 447;
                sine[105] = 448;
                sine[106] = 449;
                sine[107] = 450;
                sine[108] = 451;
                sine[109] = 452;
                sine[110] = 453;
                sine[111] = 454;
                sine[112] = 455;
                sine[113] = 456;
                sine[114] = 457;
                sine[115] = 458;
                sine[116] = 459;
                sine[117] = 460;
                sine[118] = 461;
                sine[119] = 462;
                sine[120] = 463;
                sine[121] = 464;
                sine[122] = 465;
                sine[123] = 466;
                sine[124] = 467;
                sine[125] = 468;
                sine[126] = 469;
                sine[127] = 470;
                sine[128] = 471;
                sine[129] = 472;
                sine[130] = 473;
                sine[131] = 474;
                sine[132] = 475;
                sine[133] = 476;
                sine[134] = 477;
                sine[135] = 478;
                sine[136] = 479;
                sine[137] = 480;
                sine[138] = 481;
                sine[139] = 482;
                sine[140] = 483;
                sine[141] = 483;
                sine[142] = 484;
                sine[143] = 485;
                sine[144] = 486;
                sine[145] = 487;
                sine[146] = 488;
                sine[147] = 489;
                sine[148] = 490;
                sine[149] = 491;
                sine[150] = 492;
                sine[151] = 493;
                sine[152] = 494;
                sine[153] = 495;
                sine[154] = 496;
                sine[155] = 497;
                sine[156] = 498;
                sine[157] = 498;
                sine[158] = 499;
                sine[159] = 500;
                sine[160] = 501;
                sine[161] = 502;
                sine[162] = 503;
                sine[163] = 504;
                sine[164] = 505;
                sine[165] = 506;
                sine[166] = 507;
                sine[167] = 508;
                sine[168] = 509;
                sine[169] = 509;
                sine[170] = 510;
                sine[171] = 511;
                sine[172] = 512;
                sine[173] = 513;
                sine[174] = 514;
                sine[175] = 515;
                sine[176] = 516;
                sine[177] = 517;
                sine[178] = 518;
                sine[179] = 518;
                sine[180] = 519;
                sine[181] = 520;
                sine[182] = 521;
                sine[183] = 522;
                sine[184] = 523;
                sine[185] = 524;
                sine[186] = 525;
                sine[187] = 526;
                sine[188] = 526;
                sine[189] = 527;
                sine[190] = 528;
                sine[191] = 529;
                sine[192] = 530;
                sine[193] = 531;
                sine[194] = 532;
                sine[195] = 533;
                sine[196] = 533;
                sine[197] = 534;
                sine[198] = 535;
                sine[199] = 536;
                sine[200] = 537;
                sine[201] = 538;
                sine[202] = 539;
                sine[203] = 539;
                sine[204] = 540;
                sine[205] = 541;
                sine[206] = 542;
                sine[207] = 543;
                sine[208] = 544;
                sine[209] = 544;
                sine[210] = 545;
                sine[211] = 546;
                sine[212] = 547;
                sine[213] = 548;
                sine[214] = 549;
                sine[215] = 549;
                sine[216] = 550;
                sine[217] = 551;
                sine[218] = 552;
                sine[219] = 553;
                sine[220] = 554;
                sine[221] = 554;
                sine[222] = 555;
                sine[223] = 556;
                sine[224] = 557;
                sine[225] = 558;
                sine[226] = 558;
                sine[227] = 559;
                sine[228] = 560;
                sine[229] = 561;
                sine[230] = 562;
                sine[231] = 562;
                sine[232] = 563;
                sine[233] = 564;
                sine[234] = 565;
                sine[235] = 566;
                sine[236] = 566;
                sine[237] = 567;
                sine[238] = 568;
                sine[239] = 569;
                sine[240] = 570;
                sine[241] = 570;
                sine[242] = 571;
                sine[243] = 572;
                sine[244] = 573;
                sine[245] = 573;
                sine[246] = 574;
                sine[247] = 575;
                sine[248] = 576;
                sine[249] = 576;
                sine[250] = 577;
                sine[251] = 578;
                sine[252] = 579;
                sine[253] = 579;
                sine[254] = 580;
                sine[255] = 581;
                sine[256] = 582;
                sine[257] = 582;
                sine[258] = 583;
                sine[259] = 584;
                sine[260] = 585;
                sine[261] = 585;
                sine[262] = 586;
                sine[263] = 587;
                sine[264] = 587;
                sine[265] = 588;
                sine[266] = 589;
                sine[267] = 590;
                sine[268] = 590;
                sine[269] = 591;
                sine[270] = 592;
                sine[271] = 592;
                sine[272] = 593;
                sine[273] = 594;
                sine[274] = 595;
                sine[275] = 595;
                sine[276] = 596;
                sine[277] = 597;
                sine[278] = 597;
                sine[279] = 598;
                sine[280] = 599;
                sine[281] = 599;
                sine[282] = 600;
                sine[283] = 601;
                sine[284] = 601;
                sine[285] = 602;
                sine[286] = 603;
                sine[287] = 603;
                sine[288] = 604;
                sine[289] = 605;
                sine[290] = 605;
                sine[291] = 606;
                sine[292] = 607;
                sine[293] = 607;
                sine[294] = 608;
                sine[295] = 609;
                sine[296] = 609;
                sine[297] = 610;
                sine[298] = 611;
                sine[299] = 611;
                sine[300] = 612;
                sine[301] = 613;
                sine[302] = 613;
                sine[303] = 614;
                sine[304] = 614;
                sine[305] = 615;
                sine[306] = 616;
                sine[307] = 616;
                sine[308] = 617;
                sine[309] = 617;
                sine[310] = 618;
                sine[311] = 619;
                sine[312] = 619;
                sine[313] = 620;
                sine[314] = 620;
                sine[315] = 621;
                sine[316] = 622;
                sine[317] = 622;
                sine[318] = 623;
                sine[319] = 623;
                sine[320] = 624;
                sine[321] = 625;
                sine[322] = 625;
                sine[323] = 626;
                sine[324] = 626;
                sine[325] = 627;
                sine[326] = 627;
                sine[327] = 628;
                sine[328] = 629;
                sine[329] = 629;
                sine[330] = 630;
                sine[331] = 630;
                sine[332] = 631;
                sine[333] = 631;
                sine[334] = 632;
                sine[335] = 632;
                sine[336] = 633;
                sine[337] = 634;
                sine[338] = 634;
                sine[339] = 635;
                sine[340] = 635;
                sine[341] = 636;
                sine[342] = 636;
                sine[343] = 637;
                sine[344] = 637;
                sine[345] = 638;
                sine[346] = 638;
                sine[347] = 639;
                sine[348] = 639;
                sine[349] = 640;
                sine[350] = 640;
                sine[351] = 641;
                sine[352] = 641;
                sine[353] = 642;
                sine[354] = 642;
                sine[355] = 643;
                sine[356] = 643;
                sine[357] = 644;
                sine[358] = 644;
                sine[359] = 645;
                sine[360] = 645;
                sine[361] = 646;
                sine[362] = 646;
                sine[363] = 646;
                sine[364] = 647;
                sine[365] = 647;
                sine[366] = 648;
                sine[367] = 648;
                sine[368] = 649;
                sine[369] = 649;
                sine[370] = 650;
                sine[371] = 650;
                sine[372] = 651;
                sine[373] = 651;
                sine[374] = 651;
                sine[375] = 652;
                sine[376] = 652;
                sine[377] = 653;
                sine[378] = 653;
                sine[379] = 654;
                sine[380] = 654;
                sine[381] = 654;
                sine[382] = 655;
                sine[383] = 655;
                sine[384] = 656;
                sine[385] = 656;
                sine[386] = 656;
                sine[387] = 657;
                sine[388] = 657;
                sine[389] = 658;
                sine[390] = 658;
                sine[391] = 658;
                sine[392] = 659;
                sine[393] = 659;
                sine[394] = 659;
                sine[395] = 660;
                sine[396] = 660;
                sine[397] = 660;
                sine[398] = 661;
                sine[399] = 661;
                sine[400] = 662;
                sine[401] = 662;
                sine[402] = 662;
                sine[403] = 663;
                sine[404] = 663;
                sine[405] = 663;
                sine[406] = 664;
                sine[407] = 664;
                sine[408] = 664;
                sine[409] = 665;
                sine[410] = 665;
                sine[411] = 665;
                sine[412] = 666;
                sine[413] = 666;
                sine[414] = 666;
                sine[415] = 667;
                sine[416] = 667;
                sine[417] = 667;
                sine[418] = 667;
                sine[419] = 668;
                sine[420] = 668;
                sine[421] = 668;
                sine[422] = 669;
                sine[423] = 669;
                sine[424] = 669;
                sine[425] = 669;
                sine[426] = 670;
                sine[427] = 670;
                sine[428] = 670;
                sine[429] = 671;
                sine[430] = 671;
                sine[431] = 671;
                sine[432] = 671;
                sine[433] = 672;
                sine[434] = 672;
                sine[435] = 672;
                sine[436] = 672;
                sine[437] = 673;
                sine[438] = 673;
                sine[439] = 673;
                sine[440] = 673;
                sine[441] = 673;
                sine[442] = 674;
                sine[443] = 674;
                sine[444] = 674;
                sine[445] = 674;
                sine[446] = 675;
                sine[447] = 675;
                sine[448] = 675;
                sine[449] = 675;
                sine[450] = 675;
                sine[451] = 676;
                sine[452] = 676;
                sine[453] = 676;
                sine[454] = 676;
                sine[455] = 676;
                sine[456] = 676;
                sine[457] = 677;
                sine[458] = 677;
                sine[459] = 677;
                sine[460] = 677;
                sine[461] = 677;
                sine[462] = 677;
                sine[463] = 678;
                sine[464] = 678;
                sine[465] = 678;
                sine[466] = 678;
                sine[467] = 678;
                sine[468] = 678;
                sine[469] = 679;
                sine[470] = 679;
                sine[471] = 679;
                sine[472] = 679;
                sine[473] = 679;
                sine[474] = 679;
                sine[475] = 679;
                sine[476] = 679;
                sine[477] = 680;
                sine[478] = 680;
                sine[479] = 680;
                sine[480] = 680;
                sine[481] = 680;
                sine[482] = 680;
                sine[483] = 680;
                sine[484] = 680;
                sine[485] = 680;
                sine[486] = 680;
                sine[487] = 680;
                sine[488] = 681;
                sine[489] = 681;
                sine[490] = 681;
                sine[491] = 681;
                sine[492] = 681;
                sine[493] = 681;
                sine[494] = 681;
                sine[495] = 681;
                sine[496] = 681;
                sine[497] = 681;
                sine[498] = 681;
                sine[499] = 681;
                sine[500] = 681;
                sine[501] = 681;
                sine[502] = 681;
                sine[503] = 681;
                sine[504] = 681;
                sine[505] = 681;
                sine[506] = 681;
                sine[507] = 681;
                sine[508] = 681;
                sine[509] = 681;
                sine[510] = 681;
                sine[511] = 681;
                sine[512] = 682;
                sine[513] = 681;
                sine[514] = 681;
                sine[515] = 681;
                sine[516] = 681;
                sine[517] = 681;
                sine[518] = 681;
                sine[519] = 681;
                sine[520] = 681;
                sine[521] = 681;
                sine[522] = 681;
                sine[523] = 681;
                sine[524] = 681;
                sine[525] = 681;
                sine[526] = 681;
                sine[527] = 681;
                sine[528] = 681;
                sine[529] = 681;
                sine[530] = 681;
                sine[531] = 681;
                sine[532] = 681;
                sine[533] = 681;
                sine[534] = 681;
                sine[535] = 681;
                sine[536] = 681;
                sine[537] = 680;
                sine[538] = 680;
                sine[539] = 680;
                sine[540] = 680;
                sine[541] = 680;
                sine[542] = 680;
                sine[543] = 680;
                sine[544] = 680;
                sine[545] = 680;
                sine[546] = 680;
                sine[547] = 680;
                sine[548] = 679;
                sine[549] = 679;
                sine[550] = 679;
                sine[551] = 679;
                sine[552] = 679;
                sine[553] = 679;
                sine[554] = 679;
                sine[555] = 679;
                sine[556] = 678;
                sine[557] = 678;
                sine[558] = 678;
                sine[559] = 678;
                sine[560] = 678;
                sine[561] = 678;
                sine[562] = 677;
                sine[563] = 677;
                sine[564] = 677;
                sine[565] = 677;
                sine[566] = 677;
                sine[567] = 677;
                sine[568] = 676;
                sine[569] = 676;
                sine[570] = 676;
                sine[571] = 676;
                sine[572] = 676;
                sine[573] = 676;
                sine[574] = 675;
                sine[575] = 675;
                sine[576] = 675;
                sine[577] = 675;
                sine[578] = 675;
                sine[579] = 674;
                sine[580] = 674;
                sine[581] = 674;
                sine[582] = 674;
                sine[583] = 673;
                sine[584] = 673;
                sine[585] = 673;
                sine[586] = 673;
                sine[587] = 673;
                sine[588] = 672;
                sine[589] = 672;
                sine[590] = 672;
                sine[591] = 672;
                sine[592] = 671;
                sine[593] = 671;
                sine[594] = 671;
                sine[595] = 671;
                sine[596] = 670;
                sine[597] = 670;
                sine[598] = 670;
                sine[599] = 669;
                sine[600] = 669;
                sine[601] = 669;
                sine[602] = 669;
                sine[603] = 668;
                sine[604] = 668;
                sine[605] = 668;
                sine[606] = 667;
                sine[607] = 667;
                sine[608] = 667;
                sine[609] = 667;
                sine[610] = 666;
                sine[611] = 666;
                sine[612] = 666;
                sine[613] = 665;
                sine[614] = 665;
                sine[615] = 665;
                sine[616] = 664;
                sine[617] = 664;
                sine[618] = 664;
                sine[619] = 663;
                sine[620] = 663;
                sine[621] = 663;
                sine[622] = 662;
                sine[623] = 662;
                sine[624] = 662;
                sine[625] = 661;
                sine[626] = 661;
                sine[627] = 660;
                sine[628] = 660;
                sine[629] = 660;
                sine[630] = 659;
                sine[631] = 659;
                sine[632] = 659;
                sine[633] = 658;
                sine[634] = 658;
                sine[635] = 658;
                sine[636] = 657;
                sine[637] = 657;
                sine[638] = 656;
                sine[639] = 656;
                sine[640] = 656;
                sine[641] = 655;
                sine[642] = 655;
                sine[643] = 654;
                sine[644] = 654;
                sine[645] = 654;
                sine[646] = 653;
                sine[647] = 653;
                sine[648] = 652;
                sine[649] = 652;
                sine[650] = 651;
                sine[651] = 651;
                sine[652] = 651;
                sine[653] = 650;
                sine[654] = 650;
                sine[655] = 649;
                sine[656] = 649;
                sine[657] = 648;
                sine[658] = 648;
                sine[659] = 647;
                sine[660] = 647;
                sine[661] = 646;
                sine[662] = 646;
                sine[663] = 646;
                sine[664] = 645;
                sine[665] = 645;
                sine[666] = 644;
                sine[667] = 644;
                sine[668] = 643;
                sine[669] = 643;
                sine[670] = 642;
                sine[671] = 642;
                sine[672] = 641;
                sine[673] = 641;
                sine[674] = 640;
                sine[675] = 640;
                sine[676] = 639;
                sine[677] = 639;
                sine[678] = 638;
                sine[679] = 638;
                sine[680] = 637;
                sine[681] = 637;
                sine[682] = 636;
                sine[683] = 636;
                sine[684] = 635;
                sine[685] = 635;
                sine[686] = 634;
                sine[687] = 634;
                sine[688] = 633;
                sine[689] = 632;
                sine[690] = 632;
                sine[691] = 631;
                sine[692] = 631;
                sine[693] = 630;
                sine[694] = 630;
                sine[695] = 629;
                sine[696] = 629;
                sine[697] = 628;
                sine[698] = 627;
                sine[699] = 627;
                sine[700] = 626;
                sine[701] = 626;
                sine[702] = 625;
                sine[703] = 625;
                sine[704] = 624;
                sine[705] = 623;
                sine[706] = 623;
                sine[707] = 622;
                sine[708] = 622;
                sine[709] = 621;
                sine[710] = 620;
                sine[711] = 620;
                sine[712] = 619;
                sine[713] = 619;
                sine[714] = 618;
                sine[715] = 617;
                sine[716] = 617;
                sine[717] = 616;
                sine[718] = 616;
                sine[719] = 615;
                sine[720] = 614;
                sine[721] = 614;
                sine[722] = 613;
                sine[723] = 613;
                sine[724] = 612;
                sine[725] = 611;
                sine[726] = 611;
                sine[727] = 610;
                sine[728] = 609;
                sine[729] = 609;
                sine[730] = 608;
                sine[731] = 607;
                sine[732] = 607;
                sine[733] = 606;
                sine[734] = 605;
                sine[735] = 605;
                sine[736] = 604;
                sine[737] = 603;
                sine[738] = 603;
                sine[739] = 602;
                sine[740] = 601;
                sine[741] = 601;
                sine[742] = 600;
                sine[743] = 599;
                sine[744] = 599;
                sine[745] = 598;
                sine[746] = 597;
                sine[747] = 597;
                sine[748] = 596;
                sine[749] = 595;
                sine[750] = 595;
                sine[751] = 594;
                sine[752] = 593;
                sine[753] = 592;
                sine[754] = 592;
                sine[755] = 591;
                sine[756] = 590;
                sine[757] = 590;
                sine[758] = 589;
                sine[759] = 588;
                sine[760] = 587;
                sine[761] = 587;
                sine[762] = 586;
                sine[763] = 585;
                sine[764] = 585;
                sine[765] = 584;
                sine[766] = 583;
                sine[767] = 582;
                sine[768] = 582;
                sine[769] = 581;
                sine[770] = 580;
                sine[771] = 579;
                sine[772] = 579;
                sine[773] = 578;
                sine[774] = 577;
                sine[775] = 576;
                sine[776] = 576;
                sine[777] = 575;
                sine[778] = 574;
                sine[779] = 573;
                sine[780] = 573;
                sine[781] = 572;
                sine[782] = 571;
                sine[783] = 570;
                sine[784] = 570;
                sine[785] = 569;
                sine[786] = 568;
                sine[787] = 567;
                sine[788] = 566;
                sine[789] = 566;
                sine[790] = 565;
                sine[791] = 564;
                sine[792] = 563;
                sine[793] = 562;
                sine[794] = 562;
                sine[795] = 561;
                sine[796] = 560;
                sine[797] = 559;
                sine[798] = 558;
                sine[799] = 558;
                sine[800] = 557;
                sine[801] = 556;
                sine[802] = 555;
                sine[803] = 554;
                sine[804] = 554;
                sine[805] = 553;
                sine[806] = 552;
                sine[807] = 551;
                sine[808] = 550;
                sine[809] = 549;
                sine[810] = 549;
                sine[811] = 548;
                sine[812] = 547;
                sine[813] = 546;
                sine[814] = 545;
                sine[815] = 544;
                sine[816] = 544;
                sine[817] = 543;
                sine[818] = 542;
                sine[819] = 541;
                sine[820] = 540;
                sine[821] = 539;
                sine[822] = 539;
                sine[823] = 538;
                sine[824] = 537;
                sine[825] = 536;
                sine[826] = 535;
                sine[827] = 534;
                sine[828] = 533;
                sine[829] = 533;
                sine[830] = 532;
                sine[831] = 531;
                sine[832] = 530;
                sine[833] = 529;
                sine[834] = 528;
                sine[835] = 527;
                sine[836] = 526;
                sine[837] = 526;
                sine[838] = 525;
                sine[839] = 524;
                sine[840] = 523;
                sine[841] = 522;
                sine[842] = 521;
                sine[843] = 520;
                sine[844] = 519;
                sine[845] = 518;
                sine[846] = 518;
                sine[847] = 517;
                sine[848] = 516;
                sine[849] = 515;
                sine[850] = 514;
                sine[851] = 513;
                sine[852] = 512;
                sine[853] = 511;
                sine[854] = 510;
                sine[855] = 509;
                sine[856] = 509;
                sine[857] = 508;
                sine[858] = 507;
                sine[859] = 506;
                sine[860] = 505;
                sine[861] = 504;
                sine[862] = 503;
                sine[863] = 502;
                sine[864] = 501;
                sine[865] = 500;
                sine[866] = 499;
                sine[867] = 498;
                sine[868] = 498;
                sine[869] = 497;
                sine[870] = 496;
                sine[871] = 495;
                sine[872] = 494;
                sine[873] = 493;
                sine[874] = 492;
                sine[875] = 491;
                sine[876] = 490;
                sine[877] = 489;
                sine[878] = 488;
                sine[879] = 487;
                sine[880] = 486;
                sine[881] = 485;
                sine[882] = 484;
                sine[883] = 483;
                sine[884] = 483;
                sine[885] = 482;
                sine[886] = 481;
                sine[887] = 480;
                sine[888] = 479;
                sine[889] = 478;
                sine[890] = 477;
                sine[891] = 476;
                sine[892] = 475;
                sine[893] = 474;
                sine[894] = 473;
                sine[895] = 472;
                sine[896] = 471;
                sine[897] = 470;
                sine[898] = 469;
                sine[899] = 468;
                sine[900] = 467;
                sine[901] = 466;
                sine[902] = 465;
                sine[903] = 464;
                sine[904] = 463;
                sine[905] = 462;
                sine[906] = 461;
                sine[907] = 460;
                sine[908] = 459;
                sine[909] = 458;
                sine[910] = 457;
                sine[911] = 456;
                sine[912] = 455;
                sine[913] = 454;
                sine[914] = 453;
                sine[915] = 452;
                sine[916] = 451;
                sine[917] = 450;
                sine[918] = 449;
                sine[919] = 448;
                sine[920] = 447;
                sine[921] = 446;
                sine[922] = 445;
                sine[923] = 444;
                sine[924] = 443;
                sine[925] = 442;
                sine[926] = 441;
                sine[927] = 440;
                sine[928] = 439;
                sine[929] = 438;
                sine[930] = 437;
                sine[931] = 436;
                sine[932] = 435;
                sine[933] = 434;
                sine[934] = 433;
                sine[935] = 432;
                sine[936] = 431;
                sine[937] = 430;
                sine[938] = 429;
                sine[939] = 428;
                sine[940] = 427;
                sine[941] = 426;
                sine[942] = 425;
                sine[943] = 424;
                sine[944] = 423;
                sine[945] = 422;
                sine[946] = 421;
                sine[947] = 420;
                sine[948] = 419;
                sine[949] = 418;
                sine[950] = 417;
                sine[951] = 416;
                sine[952] = 415;
                sine[953] = 414;
                sine[954] = 413;
                sine[955] = 412;
                sine[956] = 411;
                sine[957] = 410;
                sine[958] = 409;
                sine[959] = 408;
                sine[960] = 407;
                sine[961] = 406;
                sine[962] = 405;
                sine[963] = 404;
                sine[964] = 403;
                sine[965] = 402;
                sine[966] = 401;
                sine[967] = 400;
                sine[968] = 399;
                sine[969] = 398;
                sine[970] = 397;
                sine[971] = 396;
                sine[972] = 395;
                sine[973] = 394;
                sine[974] = 393;
                sine[975] = 392;
                sine[976] = 391;
                sine[977] = 390;
                sine[978] = 388;
                sine[979] = 387;
                sine[980] = 386;
                sine[981] = 385;
                sine[982] = 384;
                sine[983] = 383;
                sine[984] = 382;
                sine[985] = 381;
                sine[986] = 380;
                sine[987] = 379;
                sine[988] = 378;
                sine[989] = 377;
                sine[990] = 376;
                sine[991] = 375;
                sine[992] = 374;
                sine[993] = 373;
                sine[994] = 372;
                sine[995] = 371;
                sine[996] = 370;
                sine[997] = 369;
                sine[998] = 368;
                sine[999] = 367;
                sine[1000] = 366;
                sine[1001] = 365;
                sine[1002] = 363;
                sine[1003] = 362;
                sine[1004] = 361;
                sine[1005] = 360;
                sine[1006] = 359;
                sine[1007] = 358;
                sine[1008] = 357;
                sine[1009] = 356;
                sine[1010] = 355;
                sine[1011] = 354;
                sine[1012] = 353;
                sine[1013] = 352;
                sine[1014] = 351;
                sine[1015] = 350;
                sine[1016] = 349;
                sine[1017] = 348;
                sine[1018] = 347;
                sine[1019] = 346;
                sine[1020] = 345;
                sine[1021] = 344;
                sine[1022] = 343;
                sine[1023] = 342;
                sine[1024] = 341;
                sine[1025] = 339;
                sine[1026] = 338;
                sine[1027] = 337;
                sine[1028] = 336;
                sine[1029] = 335;
                sine[1030] = 334;
                sine[1031] = 333;
                sine[1032] = 332;
                sine[1033] = 331;
                sine[1034] = 330;
                sine[1035] = 329;
                sine[1036] = 328;
                sine[1037] = 327;
                sine[1038] = 326;
                sine[1039] = 325;
                sine[1040] = 324;
                sine[1041] = 323;
                sine[1042] = 322;
                sine[1043] = 321;
                sine[1044] = 320;
                sine[1045] = 319;
                sine[1046] = 318;
                sine[1047] = 316;
                sine[1048] = 315;
                sine[1049] = 314;
                sine[1050] = 313;
                sine[1051] = 312;
                sine[1052] = 311;
                sine[1053] = 310;
                sine[1054] = 309;
                sine[1055] = 308;
                sine[1056] = 307;
                sine[1057] = 306;
                sine[1058] = 305;
                sine[1059] = 304;
                sine[1060] = 303;
                sine[1061] = 302;
                sine[1062] = 301;
                sine[1063] = 300;
                sine[1064] = 299;
                sine[1065] = 298;
                sine[1066] = 297;
                sine[1067] = 296;
                sine[1068] = 295;
                sine[1069] = 294;
                sine[1070] = 293;
                sine[1071] = 291;
                sine[1072] = 290;
                sine[1073] = 289;
                sine[1074] = 288;
                sine[1075] = 287;
                sine[1076] = 286;
                sine[1077] = 285;
                sine[1078] = 284;
                sine[1079] = 283;
                sine[1080] = 282;
                sine[1081] = 281;
                sine[1082] = 280;
                sine[1083] = 279;
                sine[1084] = 278;
                sine[1085] = 277;
                sine[1086] = 276;
                sine[1087] = 275;
                sine[1088] = 274;
                sine[1089] = 273;
                sine[1090] = 272;
                sine[1091] = 271;
                sine[1092] = 270;
                sine[1093] = 269;
                sine[1094] = 268;
                sine[1095] = 267;
                sine[1096] = 266;
                sine[1097] = 265;
                sine[1098] = 264;
                sine[1099] = 263;
                sine[1100] = 262;
                sine[1101] = 261;
                sine[1102] = 260;
                sine[1103] = 259;
                sine[1104] = 258;
                sine[1105] = 257;
                sine[1106] = 256;
                sine[1107] = 255;
                sine[1108] = 254;
                sine[1109] = 253;
                sine[1110] = 252;
                sine[1111] = 251;
                sine[1112] = 250;
                sine[1113] = 249;
                sine[1114] = 248;
                sine[1115] = 247;
                sine[1116] = 246;
                sine[1117] = 245;
                sine[1118] = 244;
                sine[1119] = 243;
                sine[1120] = 242;
                sine[1121] = 241;
                sine[1122] = 240;
                sine[1123] = 239;
                sine[1124] = 238;
                sine[1125] = 237;
                sine[1126] = 236;
                sine[1127] = 235;
                sine[1128] = 234;
                sine[1129] = 233;
                sine[1130] = 232;
                sine[1131] = 231;
                sine[1132] = 230;
                sine[1133] = 229;
                sine[1134] = 228;
                sine[1135] = 227;
                sine[1136] = 226;
                sine[1137] = 225;
                sine[1138] = 224;
                sine[1139] = 223;
                sine[1140] = 222;
                sine[1141] = 221;
                sine[1142] = 220;
                sine[1143] = 219;
                sine[1144] = 218;
                sine[1145] = 217;
                sine[1146] = 216;
                sine[1147] = 215;
                sine[1148] = 214;
                sine[1149] = 213;
                sine[1150] = 212;
                sine[1151] = 211;
                sine[1152] = 210;
                sine[1153] = 209;
                sine[1154] = 208;
                sine[1155] = 207;
                sine[1156] = 206;
                sine[1157] = 205;
                sine[1158] = 204;
                sine[1159] = 203;
                sine[1160] = 202;
                sine[1161] = 201;
                sine[1162] = 200;
                sine[1163] = 199;
                sine[1164] = 198;
                sine[1165] = 198;
                sine[1166] = 197;
                sine[1167] = 196;
                sine[1168] = 195;
                sine[1169] = 194;
                sine[1170] = 193;
                sine[1171] = 192;
                sine[1172] = 191;
                sine[1173] = 190;
                sine[1174] = 189;
                sine[1175] = 188;
                sine[1176] = 187;
                sine[1177] = 186;
                sine[1178] = 185;
                sine[1179] = 184;
                sine[1180] = 183;
                sine[1181] = 183;
                sine[1182] = 182;
                sine[1183] = 181;
                sine[1184] = 180;
                sine[1185] = 179;
                sine[1186] = 178;
                sine[1187] = 177;
                sine[1188] = 176;
                sine[1189] = 175;
                sine[1190] = 174;
                sine[1191] = 173;
                sine[1192] = 172;
                sine[1193] = 172;
                sine[1194] = 171;
                sine[1195] = 170;
                sine[1196] = 169;
                sine[1197] = 168;
                sine[1198] = 167;
                sine[1199] = 166;
                sine[1200] = 165;
                sine[1201] = 164;
                sine[1202] = 163;
                sine[1203] = 163;
                sine[1204] = 162;
                sine[1205] = 161;
                sine[1206] = 160;
                sine[1207] = 159;
                sine[1208] = 158;
                sine[1209] = 157;
                sine[1210] = 156;
                sine[1211] = 155;
                sine[1212] = 155;
                sine[1213] = 154;
                sine[1214] = 153;
                sine[1215] = 152;
                sine[1216] = 151;
                sine[1217] = 150;
                sine[1218] = 149;
                sine[1219] = 148;
                sine[1220] = 148;
                sine[1221] = 147;
                sine[1222] = 146;
                sine[1223] = 145;
                sine[1224] = 144;
                sine[1225] = 143;
                sine[1226] = 142;
                sine[1227] = 142;
                sine[1228] = 141;
                sine[1229] = 140;
                sine[1230] = 139;
                sine[1231] = 138;
                sine[1232] = 137;
                sine[1233] = 137;
                sine[1234] = 136;
                sine[1235] = 135;
                sine[1236] = 134;
                sine[1237] = 133;
                sine[1238] = 132;
                sine[1239] = 132;
                sine[1240] = 131;
                sine[1241] = 130;
                sine[1242] = 129;
                sine[1243] = 128;
                sine[1244] = 127;
                sine[1245] = 127;
                sine[1246] = 126;
                sine[1247] = 125;
                sine[1248] = 124;
                sine[1249] = 123;
                sine[1250] = 123;
                sine[1251] = 122;
                sine[1252] = 121;
                sine[1253] = 120;
                sine[1254] = 119;
                sine[1255] = 119;
                sine[1256] = 118;
                sine[1257] = 117;
                sine[1258] = 116;
                sine[1259] = 115;
                sine[1260] = 115;
                sine[1261] = 114;
                sine[1262] = 113;
                sine[1263] = 112;
                sine[1264] = 111;
                sine[1265] = 111;
                sine[1266] = 110;
                sine[1267] = 109;
                sine[1268] = 108;
                sine[1269] = 108;
                sine[1270] = 107;
                sine[1271] = 106;
                sine[1272] = 105;
                sine[1273] = 105;
                sine[1274] = 104;
                sine[1275] = 103;
                sine[1276] = 102;
                sine[1277] = 102;
                sine[1278] = 101;
                sine[1279] = 100;
                sine[1280] = 99;
                sine[1281] = 99;
                sine[1282] = 98;
                sine[1283] = 97;
                sine[1284] = 96;
                sine[1285] = 96;
                sine[1286] = 95;
                sine[1287] = 94;
                sine[1288] = 94;
                sine[1289] = 93;
                sine[1290] = 92;
                sine[1291] = 91;
                sine[1292] = 91;
                sine[1293] = 90;
                sine[1294] = 89;
                sine[1295] = 89;
                sine[1296] = 88;
                sine[1297] = 87;
                sine[1298] = 86;
                sine[1299] = 86;
                sine[1300] = 85;
                sine[1301] = 84;
                sine[1302] = 84;
                sine[1303] = 83;
                sine[1304] = 82;
                sine[1305] = 82;
                sine[1306] = 81;
                sine[1307] = 80;
                sine[1308] = 80;
                sine[1309] = 79;
                sine[1310] = 78;
                sine[1311] = 78;
                sine[1312] = 77;
                sine[1313] = 76;
                sine[1314] = 76;
                sine[1315] = 75;
                sine[1316] = 74;
                sine[1317] = 74;
                sine[1318] = 73;
                sine[1319] = 72;
                sine[1320] = 72;
                sine[1321] = 71;
                sine[1322] = 70;
                sine[1323] = 70;
                sine[1324] = 69;
                sine[1325] = 68;
                sine[1326] = 68;
                sine[1327] = 67;
                sine[1328] = 67;
                sine[1329] = 66;
                sine[1330] = 65;
                sine[1331] = 65;
                sine[1332] = 64;
                sine[1333] = 64;
                sine[1334] = 63;
                sine[1335] = 62;
                sine[1336] = 62;
                sine[1337] = 61;
                sine[1338] = 61;
                sine[1339] = 60;
                sine[1340] = 59;
                sine[1341] = 59;
                sine[1342] = 58;
                sine[1343] = 58;
                sine[1344] = 57;
                sine[1345] = 56;
                sine[1346] = 56;
                sine[1347] = 55;
                sine[1348] = 55;
                sine[1349] = 54;
                sine[1350] = 54;
                sine[1351] = 53;
                sine[1352] = 52;
                sine[1353] = 52;
                sine[1354] = 51;
                sine[1355] = 51;
                sine[1356] = 50;
                sine[1357] = 50;
                sine[1358] = 49;
                sine[1359] = 49;
                sine[1360] = 48;
                sine[1361] = 47;
                sine[1362] = 47;
                sine[1363] = 46;
                sine[1364] = 46;
                sine[1365] = 45;
                sine[1366] = 45;
                sine[1367] = 44;
                sine[1368] = 44;
                sine[1369] = 43;
                sine[1370] = 43;
                sine[1371] = 42;
                sine[1372] = 42;
                sine[1373] = 41;
                sine[1374] = 41;
                sine[1375] = 40;
                sine[1376] = 40;
                sine[1377] = 39;
                sine[1378] = 39;
                sine[1379] = 38;
                sine[1380] = 38;
                sine[1381] = 37;
                sine[1382] = 37;
                sine[1383] = 36;
                sine[1384] = 36;
                sine[1385] = 35;
                sine[1386] = 35;
                sine[1387] = 35;
                sine[1388] = 34;
                sine[1389] = 34;
                sine[1390] = 33;
                sine[1391] = 33;
                sine[1392] = 32;
                sine[1393] = 32;
                sine[1394] = 31;
                sine[1395] = 31;
                sine[1396] = 30;
                sine[1397] = 30;
                sine[1398] = 30;
                sine[1399] = 29;
                sine[1400] = 29;
                sine[1401] = 28;
                sine[1402] = 28;
                sine[1403] = 27;
                sine[1404] = 27;
                sine[1405] = 27;
                sine[1406] = 26;
                sine[1407] = 26;
                sine[1408] = 25;
                sine[1409] = 25;
                sine[1410] = 25;
                sine[1411] = 24;
                sine[1412] = 24;
                sine[1413] = 23;
                sine[1414] = 23;
                sine[1415] = 23;
                sine[1416] = 22;
                sine[1417] = 22;
                sine[1418] = 22;
                sine[1419] = 21;
                sine[1420] = 21;
                sine[1421] = 21;
                sine[1422] = 20;
                sine[1423] = 20;
                sine[1424] = 19;
                sine[1425] = 19;
                sine[1426] = 19;
                sine[1427] = 18;
                sine[1428] = 18;
                sine[1429] = 18;
                sine[1430] = 17;
                sine[1431] = 17;
                sine[1432] = 17;
                sine[1433] = 16;
                sine[1434] = 16;
                sine[1435] = 16;
                sine[1436] = 15;
                sine[1437] = 15;
                sine[1438] = 15;
                sine[1439] = 14;
                sine[1440] = 14;
                sine[1441] = 14;
                sine[1442] = 14;
                sine[1443] = 13;
                sine[1444] = 13;
                sine[1445] = 13;
                sine[1446] = 12;
                sine[1447] = 12;
                sine[1448] = 12;
                sine[1449] = 12;
                sine[1450] = 11;
                sine[1451] = 11;
                sine[1452] = 11;
                sine[1453] = 10;
                sine[1454] = 10;
                sine[1455] = 10;
                sine[1456] = 10;
                sine[1457] = 9;
                sine[1458] = 9;
                sine[1459] = 9;
                sine[1460] = 9;
                sine[1461] = 8;
                sine[1462] = 8;
                sine[1463] = 8;
                sine[1464] = 8;
                sine[1465] = 8;
                sine[1466] = 7;
                sine[1467] = 7;
                sine[1468] = 7;
                sine[1469] = 7;
                sine[1470] = 6;
                sine[1471] = 6;
                sine[1472] = 6;
                sine[1473] = 6;
                sine[1474] = 6;
                sine[1475] = 5;
                sine[1476] = 5;
                sine[1477] = 5;
                sine[1478] = 5;
                sine[1479] = 5;
                sine[1480] = 5;
                sine[1481] = 4;
                sine[1482] = 4;
                sine[1483] = 4;
                sine[1484] = 4;
                sine[1485] = 4;
                sine[1486] = 4;
                sine[1487] = 3;
                sine[1488] = 3;
                sine[1489] = 3;
                sine[1490] = 3;
                sine[1491] = 3;
                sine[1492] = 3;
                sine[1493] = 2;
                sine[1494] = 2;
                sine[1495] = 2;
                sine[1496] = 2;
                sine[1497] = 2;
                sine[1498] = 2;
                sine[1499] = 2;
                sine[1500] = 2;
                sine[1501] = 1;
                sine[1502] = 1;
                sine[1503] = 1;
                sine[1504] = 1;
                sine[1505] = 1;
                sine[1506] = 1;
                sine[1507] = 1;
                sine[1508] = 1;
                sine[1509] = 1;
                sine[1510] = 1;
                sine[1511] = 1;
                sine[1512] = 0;
                sine[1513] = 0;
                sine[1514] = 0;
                sine[1515] = 0;
                sine[1516] = 0;
                sine[1517] = 0;
                sine[1518] = 0;
                sine[1519] = 0;
                sine[1520] = 0;
                sine[1521] = 0;
                sine[1522] = 0;
                sine[1523] = 0;
                sine[1524] = 0;
                sine[1525] = 0;
                sine[1526] = 0;
                sine[1527] = 0;
                sine[1528] = 0;
                sine[1529] = 0;
                sine[1530] = 0;
                sine[1531] = 0;
                sine[1532] = 0;
                sine[1533] = 0;
                sine[1534] = 0;
                sine[1535] = 0;
                sine[1536] = 0;
                sine[1537] = 0;
                sine[1538] = 0;
                sine[1539] = 0;
                sine[1540] = 0;
                sine[1541] = 0;
                sine[1542] = 0;
                sine[1543] = 0;
                sine[1544] = 0;
                sine[1545] = 0;
                sine[1546] = 0;
                sine[1547] = 0;
                sine[1548] = 0;
                sine[1549] = 0;
                sine[1550] = 0;
                sine[1551] = 0;
                sine[1552] = 0;
                sine[1553] = 0;
                sine[1554] = 0;
                sine[1555] = 0;
                sine[1556] = 0;
                sine[1557] = 0;
                sine[1558] = 0;
                sine[1559] = 0;
                sine[1560] = 0;
                sine[1561] = 1;
                sine[1562] = 1;
                sine[1563] = 1;
                sine[1564] = 1;
                sine[1565] = 1;
                sine[1566] = 1;
                sine[1567] = 1;
                sine[1568] = 1;
                sine[1569] = 1;
                sine[1570] = 1;
                sine[1571] = 1;
                sine[1572] = 2;
                sine[1573] = 2;
                sine[1574] = 2;
                sine[1575] = 2;
                sine[1576] = 2;
                sine[1577] = 2;
                sine[1578] = 2;
                sine[1579] = 2;
                sine[1580] = 3;
                sine[1581] = 3;
                sine[1582] = 3;
                sine[1583] = 3;
                sine[1584] = 3;
                sine[1585] = 3;
                sine[1586] = 4;
                sine[1587] = 4;
                sine[1588] = 4;
                sine[1589] = 4;
                sine[1590] = 4;
                sine[1591] = 4;
                sine[1592] = 5;
                sine[1593] = 5;
                sine[1594] = 5;
                sine[1595] = 5;
                sine[1596] = 5;
                sine[1597] = 5;
                sine[1598] = 6;
                sine[1599] = 6;
                sine[1600] = 6;
                sine[1601] = 6;
                sine[1602] = 6;
                sine[1603] = 7;
                sine[1604] = 7;
                sine[1605] = 7;
                sine[1606] = 7;
                sine[1607] = 8;
                sine[1608] = 8;
                sine[1609] = 8;
                sine[1610] = 8;
                sine[1611] = 8;
                sine[1612] = 9;
                sine[1613] = 9;
                sine[1614] = 9;
                sine[1615] = 9;
                sine[1616] = 10;
                sine[1617] = 10;
                sine[1618] = 10;
                sine[1619] = 10;
                sine[1620] = 11;
                sine[1621] = 11;
                sine[1622] = 11;
                sine[1623] = 12;
                sine[1624] = 12;
                sine[1625] = 12;
                sine[1626] = 12;
                sine[1627] = 13;
                sine[1628] = 13;
                sine[1629] = 13;
                sine[1630] = 14;
                sine[1631] = 14;
                sine[1632] = 14;
                sine[1633] = 14;
                sine[1634] = 15;
                sine[1635] = 15;
                sine[1636] = 15;
                sine[1637] = 16;
                sine[1638] = 16;
                sine[1639] = 16;
                sine[1640] = 17;
                sine[1641] = 17;
                sine[1642] = 17;
                sine[1643] = 18;
                sine[1644] = 18;
                sine[1645] = 18;
                sine[1646] = 19;
                sine[1647] = 19;
                sine[1648] = 19;
                sine[1649] = 20;
                sine[1650] = 20;
                sine[1651] = 21;
                sine[1652] = 21;
                sine[1653] = 21;
                sine[1654] = 22;
                sine[1655] = 22;
                sine[1656] = 22;
                sine[1657] = 23;
                sine[1658] = 23;
                sine[1659] = 23;
                sine[1660] = 24;
                sine[1661] = 24;
                sine[1662] = 25;
                sine[1663] = 25;
                sine[1664] = 25;
                sine[1665] = 26;
                sine[1666] = 26;
                sine[1667] = 27;
                sine[1668] = 27;
                sine[1669] = 27;
                sine[1670] = 28;
                sine[1671] = 28;
                sine[1672] = 29;
                sine[1673] = 29;
                sine[1674] = 30;
                sine[1675] = 30;
                sine[1676] = 30;
                sine[1677] = 31;
                sine[1678] = 31;
                sine[1679] = 32;
                sine[1680] = 32;
                sine[1681] = 33;
                sine[1682] = 33;
                sine[1683] = 34;
                sine[1684] = 34;
                sine[1685] = 35;
                sine[1686] = 35;
                sine[1687] = 35;
                sine[1688] = 36;
                sine[1689] = 36;
                sine[1690] = 37;
                sine[1691] = 37;
                sine[1692] = 38;
                sine[1693] = 38;
                sine[1694] = 39;
                sine[1695] = 39;
                sine[1696] = 40;
                sine[1697] = 40;
                sine[1698] = 41;
                sine[1699] = 41;
                sine[1700] = 42;
                sine[1701] = 42;
                sine[1702] = 43;
                sine[1703] = 43;
                sine[1704] = 44;
                sine[1705] = 44;
                sine[1706] = 45;
                sine[1707] = 45;
                sine[1708] = 46;
                sine[1709] = 46;
                sine[1710] = 47;
                sine[1711] = 47;
                sine[1712] = 48;
                sine[1713] = 49;
                sine[1714] = 49;
                sine[1715] = 50;
                sine[1716] = 50;
                sine[1717] = 51;
                sine[1718] = 51;
                sine[1719] = 52;
                sine[1720] = 52;
                sine[1721] = 53;
                sine[1722] = 54;
                sine[1723] = 54;
                sine[1724] = 55;
                sine[1725] = 55;
                sine[1726] = 56;
                sine[1727] = 56;
                sine[1728] = 57;
                sine[1729] = 58;
                sine[1730] = 58;
                sine[1731] = 59;
                sine[1732] = 59;
                sine[1733] = 60;
                sine[1734] = 61;
                sine[1735] = 61;
                sine[1736] = 62;
                sine[1737] = 62;
                sine[1738] = 63;
                sine[1739] = 64;
                sine[1740] = 64;
                sine[1741] = 65;
                sine[1742] = 65;
                sine[1743] = 66;
                sine[1744] = 67;
                sine[1745] = 67;
                sine[1746] = 68;
                sine[1747] = 68;
                sine[1748] = 69;
                sine[1749] = 70;
                sine[1750] = 70;
                sine[1751] = 71;
                sine[1752] = 72;
                sine[1753] = 72;
                sine[1754] = 73;
                sine[1755] = 74;
                sine[1756] = 74;
                sine[1757] = 75;
                sine[1758] = 76;
                sine[1759] = 76;
                sine[1760] = 77;
                sine[1761] = 78;
                sine[1762] = 78;
                sine[1763] = 79;
                sine[1764] = 80;
                sine[1765] = 80;
                sine[1766] = 81;
                sine[1767] = 82;
                sine[1768] = 82;
                sine[1769] = 83;
                sine[1770] = 84;
                sine[1771] = 84;
                sine[1772] = 85;
                sine[1773] = 86;
                sine[1774] = 86;
                sine[1775] = 87;
                sine[1776] = 88;
                sine[1777] = 89;
                sine[1778] = 89;
                sine[1779] = 90;
                sine[1780] = 91;
                sine[1781] = 91;
                sine[1782] = 92;
                sine[1783] = 93;
                sine[1784] = 94;
                sine[1785] = 94;
                sine[1786] = 95;
                sine[1787] = 96;
                sine[1788] = 96;
                sine[1789] = 97;
                sine[1790] = 98;
                sine[1791] = 99;
                sine[1792] = 99;
                sine[1793] = 100;
                sine[1794] = 101;
                sine[1795] = 102;
                sine[1796] = 102;
                sine[1797] = 103;
                sine[1798] = 104;
                sine[1799] = 105;
                sine[1800] = 105;
                sine[1801] = 106;
                sine[1802] = 107;
                sine[1803] = 108;
                sine[1804] = 108;
                sine[1805] = 109;
                sine[1806] = 110;
                sine[1807] = 111;
                sine[1808] = 111;
                sine[1809] = 112;
                sine[1810] = 113;
                sine[1811] = 114;
                sine[1812] = 115;
                sine[1813] = 115;
                sine[1814] = 116;
                sine[1815] = 117;
                sine[1816] = 118;
                sine[1817] = 119;
                sine[1818] = 119;
                sine[1819] = 120;
                sine[1820] = 121;
                sine[1821] = 122;
                sine[1822] = 123;
                sine[1823] = 123;
                sine[1824] = 124;
                sine[1825] = 125;
                sine[1826] = 126;
                sine[1827] = 127;
                sine[1828] = 127;
                sine[1829] = 128;
                sine[1830] = 129;
                sine[1831] = 130;
                sine[1832] = 131;
                sine[1833] = 132;
                sine[1834] = 132;
                sine[1835] = 133;
                sine[1836] = 134;
                sine[1837] = 135;
                sine[1838] = 136;
                sine[1839] = 137;
                sine[1840] = 137;
                sine[1841] = 138;
                sine[1842] = 139;
                sine[1843] = 140;
                sine[1844] = 141;
                sine[1845] = 142;
                sine[1846] = 142;
                sine[1847] = 143;
                sine[1848] = 144;
                sine[1849] = 145;
                sine[1850] = 146;
                sine[1851] = 147;
                sine[1852] = 148;
                sine[1853] = 148;
                sine[1854] = 149;
                sine[1855] = 150;
                sine[1856] = 151;
                sine[1857] = 152;
                sine[1858] = 153;
                sine[1859] = 154;
                sine[1860] = 155;
                sine[1861] = 155;
                sine[1862] = 156;
                sine[1863] = 157;
                sine[1864] = 158;
                sine[1865] = 159;
                sine[1866] = 160;
                sine[1867] = 161;
                sine[1868] = 162;
                sine[1869] = 163;
                sine[1870] = 163;
                sine[1871] = 164;
                sine[1872] = 165;
                sine[1873] = 166;
                sine[1874] = 167;
                sine[1875] = 168;
                sine[1876] = 169;
                sine[1877] = 170;
                sine[1878] = 171;
                sine[1879] = 172;
                sine[1880] = 172;
                sine[1881] = 173;
                sine[1882] = 174;
                sine[1883] = 175;
                sine[1884] = 176;
                sine[1885] = 177;
                sine[1886] = 178;
                sine[1887] = 179;
                sine[1888] = 180;
                sine[1889] = 181;
                sine[1890] = 182;
                sine[1891] = 183;
                sine[1892] = 183;
                sine[1893] = 184;
                sine[1894] = 185;
                sine[1895] = 186;
                sine[1896] = 187;
                sine[1897] = 188;
                sine[1898] = 189;
                sine[1899] = 190;
                sine[1900] = 191;
                sine[1901] = 192;
                sine[1902] = 193;
                sine[1903] = 194;
                sine[1904] = 195;
                sine[1905] = 196;
                sine[1906] = 197;
                sine[1907] = 198;
                sine[1908] = 198;
                sine[1909] = 199;
                sine[1910] = 200;
                sine[1911] = 201;
                sine[1912] = 202;
                sine[1913] = 203;
                sine[1914] = 204;
                sine[1915] = 205;
                sine[1916] = 206;
                sine[1917] = 207;
                sine[1918] = 208;
                sine[1919] = 209;
                sine[1920] = 210;
                sine[1921] = 211;
                sine[1922] = 212;
                sine[1923] = 213;
                sine[1924] = 214;
                sine[1925] = 215;
                sine[1926] = 216;
                sine[1927] = 217;
                sine[1928] = 218;
                sine[1929] = 219;
                sine[1930] = 220;
                sine[1931] = 221;
                sine[1932] = 222;
                sine[1933] = 223;
                sine[1934] = 224;
                sine[1935] = 225;
                sine[1936] = 226;
                sine[1937] = 227;
                sine[1938] = 228;
                sine[1939] = 229;
                sine[1940] = 230;
                sine[1941] = 231;
                sine[1942] = 232;
                sine[1943] = 233;
                sine[1944] = 234;
                sine[1945] = 235;
                sine[1946] = 236;
                sine[1947] = 237;
                sine[1948] = 238;
                sine[1949] = 239;
                sine[1950] = 240;
                sine[1951] = 241;
                sine[1952] = 242;
                sine[1953] = 243;
                sine[1954] = 244;
                sine[1955] = 245;
                sine[1956] = 246;
                sine[1957] = 247;
                sine[1958] = 248;
                sine[1959] = 249;
                sine[1960] = 250;
                sine[1961] = 251;
                sine[1962] = 252;
                sine[1963] = 253;
                sine[1964] = 254;
                sine[1965] = 255;
                sine[1966] = 256;
                sine[1967] = 257;
                sine[1968] = 258;
                sine[1969] = 259;
                sine[1970] = 260;
                sine[1971] = 261;
                sine[1972] = 262;
                sine[1973] = 263;
                sine[1974] = 264;
                sine[1975] = 265;
                sine[1976] = 266;
                sine[1977] = 267;
                sine[1978] = 268;
                sine[1979] = 269;
                sine[1980] = 270;
                sine[1981] = 271;
                sine[1982] = 272;
                sine[1983] = 273;
                sine[1984] = 274;
                sine[1985] = 275;
                sine[1986] = 276;
                sine[1987] = 277;
                sine[1988] = 278;
                sine[1989] = 279;
                sine[1990] = 280;
                sine[1991] = 281;
                sine[1992] = 282;
                sine[1993] = 283;
                sine[1994] = 284;
                sine[1995] = 285;
                sine[1996] = 286;
                sine[1997] = 287;
                sine[1998] = 288;
                sine[1999] = 289;
                sine[2000] = 290;
                sine[2001] = 291;
                sine[2002] = 293;
                sine[2003] = 294;
                sine[2004] = 295;
                sine[2005] = 296;
                sine[2006] = 297;
                sine[2007] = 298;
                sine[2008] = 299;
                sine[2009] = 300;
                sine[2010] = 301;
                sine[2011] = 302;
                sine[2012] = 303;
                sine[2013] = 304;
                sine[2014] = 305;
                sine[2015] = 306;
                sine[2016] = 307;
                sine[2017] = 308;
                sine[2018] = 309;
                sine[2019] = 310;
                sine[2020] = 311;
                sine[2021] = 312;
                sine[2022] = 313;
                sine[2023] = 314;
                sine[2024] = 315;
                sine[2025] = 316;
                sine[2026] = 318;
                sine[2027] = 319;
                sine[2028] = 320;
                sine[2029] = 321;
                sine[2030] = 322;
                sine[2031] = 323;
                sine[2032] = 324;
                sine[2033] = 325;
                sine[2034] = 326;
                sine[2035] = 327;
                sine[2036] = 328;
                sine[2037] = 329;
                sine[2038] = 330;
                sine[2039] = 331;
                sine[2040] = 332;
                sine[2041] = 333;
                sine[2042] = 334;
                sine[2043] = 335;
                sine[2044] = 336;
                sine[2045] = 337;
                sine[2046] = 338;
                sine[2047] = 339;   
    end
endmodule
